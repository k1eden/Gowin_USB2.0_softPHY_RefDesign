`timescale 100 ps/100 ps
module USB_Device_Controller_Top (
  clk_i,
  reset_i,
  usbrst_o,
  highspeed_o,
  suspend_o,
  online_o,
  txdat_i,
  txval_i,
  txdat_len_i,
  txiso_pid_i,
  txcork_i,
  txpop_o,
  txact_o,
  txpktfin_o,
  rxdat_o,
  rxval_o,
  rxrdy_i,
  rxact_o,
  rxpktval_o,
  setup_o,
  endpt_o,
  sof_o,
  inf_alter_i,
  inf_alter_o,
  inf_sel_o,
  inf_set_o,
  descrom_raddr_o,
  descrom_rdata_i,
  desc_dev_addr_i,
  desc_dev_len_i,
  desc_qual_addr_i,
  desc_qual_len_i,
  desc_fscfg_addr_i,
  desc_fscfg_len_i,
  desc_hscfg_addr_i,
  desc_hscfg_len_i,
  desc_oscfg_addr_i,
  desc_strlang_addr_i,
  desc_strvendor_addr_i,
  desc_strvendor_len_i,
  desc_strproduct_addr_i,
  desc_strproduct_len_i,
  desc_strserial_addr_i,
  desc_strserial_len_i,
  desc_have_strings_i,
  utmi_dataout_o,
  utmi_txvalid_o,
  utmi_txready_i,
  utmi_datain_i,
  utmi_rxactive_i,
  utmi_rxvalid_i,
  utmi_rxerror_i,
  utmi_linestate_i,
  utmi_opmode_o,
  utmi_xcvrselect_o,
  utmi_termselect_o,
  utmi_reset_o
)
;
input clk_i;
input reset_i;
output usbrst_o;
output highspeed_o;
output suspend_o;
output online_o;
input [7:0] txdat_i;
input txval_i;
input [11:0] txdat_len_i;
input [3:0] txiso_pid_i;
input txcork_i;
output txpop_o;
output txact_o;
output txpktfin_o;
output [7:0] rxdat_o;
output rxval_o;
input rxrdy_i;
output rxact_o;
output rxpktval_o;
output setup_o;
output [3:0] endpt_o;
output sof_o;
input [7:0] inf_alter_i;
output [7:0] inf_alter_o;
output [7:0] inf_sel_o;
output inf_set_o;
output [9:0] descrom_raddr_o;
input [7:0] descrom_rdata_i;
input [9:0] desc_dev_addr_i;
input [7:0] desc_dev_len_i;
input [9:0] desc_qual_addr_i;
input [7:0] desc_qual_len_i;
input [9:0] desc_fscfg_addr_i;
input [7:0] desc_fscfg_len_i;
input [9:0] desc_hscfg_addr_i;
input [7:0] desc_hscfg_len_i;
input [9:0] desc_oscfg_addr_i;
input [9:0] desc_strlang_addr_i;
input [9:0] desc_strvendor_addr_i;
input [7:0] desc_strvendor_len_i;
input [9:0] desc_strproduct_addr_i;
input [7:0] desc_strproduct_len_i;
input [9:0] desc_strserial_addr_i;
input [7:0] desc_strserial_len_i;
input desc_have_strings_i;
output [7:0] utmi_dataout_o;
output utmi_txvalid_o;
input utmi_txready_i;
input [7:0] utmi_datain_i;
input utmi_rxactive_i;
input utmi_rxvalid_i;
input utmi_rxerror_i;
input [1:0] utmi_linestate_i;
output [1:0] utmi_opmode_o;
output [1:0] utmi_xcvrselect_o;
output utmi_termselect_o;
output utmi_reset_o;
wire clk_i_d;
wire reset_i_d;
wire txval_i_d;
wire txcork_i_d;
wire rxrdy_i_d;
wire desc_have_strings_i_d;
wire utmi_txready_i_d;
wire utmi_rxactive_i_d;
wire utmi_rxvalid_i_d;
wire utmi_rxerror_i_d;
wire u_usb_device_controller_usb_transact_inst_T_PING_2;
wire u_usb_device_controller_usb_transact_inst_s_setup_2;
wire u_usb_device_controller_s_endpt_rxrdy;
wire u_usb_device_controller_s_endpt_txcork;
wire u_usb_device_controller_s_halt_out;
wire u_usb_device_controller_s_halt_in;
wire u_usb_device_controller_s_osync;
wire u_usb_device_controller_s_isync;
wire u_usb_device_controller_rxval_d2;
wire u_usb_device_controller_rxpktval_o_d;
wire u_usb_device_controller_test_packet_inst_test_en_dly_Z;
wire u_usb_device_controller_test_packet_inst_test_en_dect;
wire u_usb_device_controller_u_usb_init_v_clrtimer2;
wire u_usb_device_controller_u_usb_init_utmi_reset_o_d;
wire u_usb_device_controller_u_usb_init_usbp_chirpk;
wire u_usb_device_controller_u_usb_init_highspeed_o_d;
wire u_usb_device_controller_u_usb_init_suspend_o_d;
wire u_usb_device_controller_u_usb_init_v_clrtimer1;
wire u_usb_device_controller_u_usb_packet_s_txfirst;
wire u_usb_device_controller_u_usb_packet_usbp_rxact;
wire u_usb_device_controller_u_usb_packet_s_rxvalid;
wire u_usb_device_controller_u_usb_packet_s_rxerror;
wire u_usb_device_controller_u_usb_packet_s_txready;
wire u_usb_device_controller_u_usb_packet_s_rxgoodpacket;
wire u_usb_device_controller_usb_transact_inst_s_setup;
wire u_usb_device_controller_usb_transact_inst_usbt_osync;
wire u_usb_device_controller_usb_transact_inst_s_prevrxact;
wire u_usb_device_controller_usb_control_inst_online_o_d;
wire u_usb_device_controller_usb_control_inst_usbc_test_en;
wire u_usb_device_controller_usb_control_inst_s_test_sel;
wire u_usb_device_controller_rxval_d0;
wire u_usb_device_controller_rxval_d1;
wire u_usb_device_controller_u_usb_init_utmi_termselect_o_d;
wire u_usb_device_controller_u_usb_packet_usbp_txvalid_o;
wire u_usb_device_controller_txact_o_d;
wire u_usb_device_controller_s_nyet;
wire u_usb_device_controller_usb_transact_inst_s_in;
wire u_usb_device_controller_usb_transact_inst_s_out;
wire u_usb_device_controller_usb_transact_inst_s_sof;
wire u_usb_device_controller_usb_transact_inst_s_in_valid;
wire u_usb_device_controller_usb_transact_inst_s_out_valid;
wire u_usb_device_controller_usb_transact_inst_sof_o_d;
wire u_usb_device_controller_usb_transact_inst_s_ping;
wire u_usb_device_controller_usb_transact_inst_usbt_fin;
wire u_usb_device_controller_usb_control_inst_inf_set_o_d;
wire u_usb_device_controller_n1473;
wire u_usb_device_controller_n1473_28;
wire u_usb_device_controller_n1473_29;
wire u_usb_device_controller_n1473_30;
wire u_usb_device_controller_n1473_31;
wire u_usb_device_controller_n1473_32;
wire u_usb_device_controller_n1473_33;
wire u_usb_device_controller_n1473_34;
wire u_usb_device_controller_n1473_35;
wire u_usb_device_controller_n1473_36;
wire u_usb_device_controller_n1473_37;
wire u_usb_device_controller_n1473_38;
wire u_usb_device_controller_n1473_39;
wire u_usb_device_controller_n1473_40;
wire u_usb_device_controller_n1473_41;
wire u_usb_device_controller_n1473_42;
wire u_usb_device_controller_n1473_43;
wire u_usb_device_controller_n1473_44;
wire u_usb_device_controller_n1473_45;
wire u_usb_device_controller_n1473_46;
wire u_usb_device_controller_n1473_47;
wire u_usb_device_controller_n1473_48;
wire u_usb_device_controller_n1473_49;
wire u_usb_device_controller_n1473_50;
wire u_usb_device_controller_n2023;
wire u_usb_device_controller_n2023_2;
wire u_usb_device_controller_n2022;
wire u_usb_device_controller_n2022_2;
wire u_usb_device_controller_n2021;
wire u_usb_device_controller_n2021_2;
wire u_usb_device_controller_n2020;
wire u_usb_device_controller_n2020_2;
wire u_usb_device_controller_n2019;
wire u_usb_device_controller_n2019_2;
wire u_usb_device_controller_n2018;
wire u_usb_device_controller_n2018_2;
wire u_usb_device_controller_n2017;
wire u_usb_device_controller_n2017_2;
wire u_usb_device_controller_n2016;
wire u_usb_device_controller_n2016_2;
wire u_usb_device_controller_n2015;
wire u_usb_device_controller_n2015_2;
wire u_usb_device_controller_u_usb_init_n240;
wire u_usb_device_controller_u_usb_init_n240_2;
wire u_usb_device_controller_u_usb_init_n239;
wire u_usb_device_controller_u_usb_init_n239_2;
wire u_usb_device_controller_u_usb_init_n238;
wire u_usb_device_controller_u_usb_init_n238_2;
wire u_usb_device_controller_u_usb_init_n237;
wire u_usb_device_controller_u_usb_init_n237_2;
wire u_usb_device_controller_u_usb_init_n236;
wire u_usb_device_controller_u_usb_init_n236_2;
wire u_usb_device_controller_u_usb_init_n235;
wire u_usb_device_controller_u_usb_init_n235_2;
wire u_usb_device_controller_u_usb_init_n234;
wire u_usb_device_controller_u_usb_init_n234_2;
wire u_usb_device_controller_u_usb_init_n233;
wire u_usb_device_controller_u_usb_init_n233_2;
wire u_usb_device_controller_u_usb_init_n232;
wire u_usb_device_controller_u_usb_init_n232_2;
wire u_usb_device_controller_u_usb_init_n231;
wire u_usb_device_controller_u_usb_init_n231_2;
wire u_usb_device_controller_u_usb_init_n230;
wire u_usb_device_controller_u_usb_init_n230_2;
wire u_usb_device_controller_u_usb_init_n229;
wire u_usb_device_controller_u_usb_init_n229_2;
wire u_usb_device_controller_u_usb_init_n228;
wire u_usb_device_controller_u_usb_init_n228_2;
wire u_usb_device_controller_u_usb_init_n227;
wire u_usb_device_controller_u_usb_init_n227_2;
wire u_usb_device_controller_u_usb_init_n226;
wire u_usb_device_controller_u_usb_init_n226_2;
wire u_usb_device_controller_u_usb_init_n278;
wire u_usb_device_controller_u_usb_init_n278_2;
wire u_usb_device_controller_u_usb_init_n277;
wire u_usb_device_controller_u_usb_init_n277_2;
wire u_usb_device_controller_u_usb_init_n276;
wire u_usb_device_controller_u_usb_init_n276_2;
wire u_usb_device_controller_u_usb_init_n275;
wire u_usb_device_controller_u_usb_init_n275_2;
wire u_usb_device_controller_u_usb_init_n274;
wire u_usb_device_controller_u_usb_init_n274_2;
wire u_usb_device_controller_u_usb_init_n273;
wire u_usb_device_controller_u_usb_init_n273_2;
wire u_usb_device_controller_u_usb_init_n272;
wire u_usb_device_controller_u_usb_init_n272_2;
wire u_usb_device_controller_u_usb_init_n271;
wire u_usb_device_controller_u_usb_init_n271_2;
wire u_usb_device_controller_u_usb_init_n270;
wire u_usb_device_controller_u_usb_init_n270_2;
wire u_usb_device_controller_u_usb_init_n269;
wire u_usb_device_controller_u_usb_init_n269_2;
wire u_usb_device_controller_u_usb_init_n268;
wire u_usb_device_controller_u_usb_init_n268_2;
wire u_usb_device_controller_u_usb_init_n267;
wire u_usb_device_controller_u_usb_init_n267_2;
wire u_usb_device_controller_u_usb_init_n266;
wire u_usb_device_controller_u_usb_init_n266_2;
wire u_usb_device_controller_u_usb_init_n265;
wire u_usb_device_controller_u_usb_init_n265_2;
wire u_usb_device_controller_u_usb_init_n264;
wire u_usb_device_controller_u_usb_init_n264_2;
wire u_usb_device_controller_u_usb_init_n263;
wire u_usb_device_controller_u_usb_init_n263_2;
wire u_usb_device_controller_u_usb_init_n262;
wire u_usb_device_controller_u_usb_init_n262_2;
wire u_usb_device_controller_u_usb_init_n261;
wire u_usb_device_controller_u_usb_init_n261_2;
wire u_usb_device_controller_u_usb_init_n260;
wire u_usb_device_controller_u_usb_init_n260_2;
wire u_usb_device_controller_test_packet_inst_test_dval;
wire u_usb_device_controller_u_usb_init_s_state_0_4;
wire u_usb_device_controller_n1454;
wire u_usb_device_controller_n1454_3;
wire u_usb_device_controller_n1455;
wire u_usb_device_controller_n1455_3;
wire u_usb_device_controller_n1456;
wire u_usb_device_controller_n1456_3;
wire u_usb_device_controller_n1457;
wire u_usb_device_controller_n1457_3;
wire u_usb_device_controller_n1458;
wire u_usb_device_controller_n1458_3;
wire u_usb_device_controller_n1459;
wire u_usb_device_controller_n1459_3;
wire u_usb_device_controller_n1460;
wire u_usb_device_controller_n1460_3;
wire u_usb_device_controller_n1461;
wire u_usb_device_controller_n1461_3;
wire u_usb_device_controller_n1462;
wire u_usb_device_controller_n1462_3;
wire u_usb_device_controller_n1463;
wire u_usb_device_controller_n1463_3;
wire u_usb_device_controller_n1464;
wire u_usb_device_controller_n1464_3;
wire u_usb_device_controller_n1465;
wire u_usb_device_controller_n1465_3;
wire u_usb_device_controller_usb_transact_inst_n156;
wire u_usb_device_controller_usb_transact_inst_n156_3;
wire u_usb_device_controller_usb_transact_inst_n157;
wire u_usb_device_controller_usb_transact_inst_n157_3;
wire u_usb_device_controller_usb_transact_inst_n158;
wire u_usb_device_controller_usb_transact_inst_n158_3;
wire u_usb_device_controller_usb_transact_inst_n159;
wire u_usb_device_controller_usb_transact_inst_n159_3;
wire u_usb_device_controller_usb_transact_inst_n160;
wire u_usb_device_controller_usb_transact_inst_n160_3;
wire u_usb_device_controller_usb_transact_inst_n161;
wire u_usb_device_controller_usb_transact_inst_n161_3;
wire u_usb_device_controller_usb_transact_inst_n162;
wire u_usb_device_controller_usb_transact_inst_n162_3;
wire u_usb_device_controller_usb_control_inst_n1467;
wire u_usb_device_controller_usb_control_inst_n1467_3;
wire u_usb_device_controller_usb_control_inst_n1468;
wire u_usb_device_controller_usb_control_inst_n1468_3;
wire u_usb_device_controller_usb_control_inst_n1469;
wire u_usb_device_controller_usb_control_inst_n1469_3;
wire u_usb_device_controller_usb_control_inst_n1470;
wire u_usb_device_controller_usb_control_inst_n1470_3;
wire u_usb_device_controller_usb_control_inst_n1471;
wire u_usb_device_controller_usb_control_inst_n1471_3;
wire u_usb_device_controller_usb_control_inst_n1472;
wire u_usb_device_controller_usb_control_inst_n1472_3;
wire u_usb_device_controller_usb_control_inst_n1473;
wire u_usb_device_controller_usb_control_inst_n1473_3;
wire u_usb_device_controller_usb_control_inst_n1474;
wire u_usb_device_controller_usb_control_inst_n1474_3;
wire u_usb_device_controller_usb_control_inst_n1476;
wire u_usb_device_controller_usb_control_inst_n1476_3;
wire u_usb_device_controller_usb_control_inst_n1477;
wire u_usb_device_controller_usb_control_inst_n1477_3;
wire u_usb_device_controller_usb_control_inst_n1478;
wire u_usb_device_controller_usb_control_inst_n1478_3;
wire u_usb_device_controller_usb_control_inst_n1479;
wire u_usb_device_controller_usb_control_inst_n1479_3;
wire u_usb_device_controller_usb_control_inst_n1480;
wire u_usb_device_controller_usb_control_inst_n1480_3;
wire u_usb_device_controller_usb_control_inst_n1481;
wire u_usb_device_controller_usb_control_inst_n1481_3;
wire u_usb_device_controller_usb_control_inst_n1482;
wire u_usb_device_controller_usb_control_inst_n1482_3;
wire u_usb_device_controller_usb_control_inst_n1483;
wire u_usb_device_controller_usb_control_inst_n1483_3;
wire u_usb_device_controller_usb_control_inst_n611;
wire u_usb_device_controller_usb_control_inst_n613;
wire u_usb_device_controller_usb_control_inst_n615;
wire u_usb_device_controller_usb_control_inst_n617;
wire u_usb_device_controller_usb_control_inst_n619;
wire u_usb_device_controller_usb_control_inst_n621;
wire u_usb_device_controller_usb_control_inst_n623;
wire u_usb_device_controller_usb_control_inst_n625;
wire u_usb_device_controller_usb_control_inst_n627;
wire u_usb_device_controller_usb_control_inst_n629;
wire u_usb_device_controller_usb_control_inst_n631;
wire u_usb_device_controller_usb_control_inst_n633;
wire u_usb_device_controller_usb_control_inst_n635;
wire u_usb_device_controller_usb_control_inst_n637;
wire u_usb_device_controller_n1241_39;
wire u_usb_device_controller_n1241_40;
wire u_usb_device_controller_n1241_41;
wire u_usb_device_controller_n1241_42;
wire u_usb_device_controller_n1241_43;
wire u_usb_device_controller_n1241_44;
wire u_usb_device_controller_n1242_39;
wire u_usb_device_controller_n1242_40;
wire u_usb_device_controller_n1242_41;
wire u_usb_device_controller_n1242_42;
wire u_usb_device_controller_n1242_43;
wire u_usb_device_controller_n1242_44;
wire u_usb_device_controller_n1243_39;
wire u_usb_device_controller_n1243_40;
wire u_usb_device_controller_n1243_41;
wire u_usb_device_controller_n1243_42;
wire u_usb_device_controller_n1243_43;
wire u_usb_device_controller_n1243_44;
wire u_usb_device_controller_n1244_39;
wire u_usb_device_controller_n1244_40;
wire u_usb_device_controller_n1244_41;
wire u_usb_device_controller_n1244_42;
wire u_usb_device_controller_n1244_43;
wire u_usb_device_controller_n1244_44;
wire u_usb_device_controller_usb_control_inst_n645;
wire u_usb_device_controller_usb_control_inst_n645_33;
wire u_usb_device_controller_usb_control_inst_n645_35;
wire u_usb_device_controller_usb_control_inst_n645_37;
wire u_usb_device_controller_usb_control_inst_n645_39;
wire u_usb_device_controller_usb_control_inst_n645_41;
wire u_usb_device_controller_usb_control_inst_n645_43;
wire u_usb_device_controller_n1241_46;
wire u_usb_device_controller_n1241_48;
wire u_usb_device_controller_n1241_50;
wire u_usb_device_controller_n1242_46;
wire u_usb_device_controller_n1242_48;
wire u_usb_device_controller_n1242_50;
wire u_usb_device_controller_n1243_46;
wire u_usb_device_controller_n1243_48;
wire u_usb_device_controller_n1243_50;
wire u_usb_device_controller_n1244_46;
wire u_usb_device_controller_n1244_48;
wire u_usb_device_controller_n1244_50;
wire u_usb_device_controller_n1241_52;
wire u_usb_device_controller_n1242_52;
wire u_usb_device_controller_n1243_52;
wire u_usb_device_controller_n1244_52;
wire u_usb_device_controller_usb_control_inst_n645_45;
wire u_usb_device_controller_usb_control_inst_n645_47;
wire u_usb_device_controller_usb_control_inst_n645_49;
wire u_usb_device_controller_usb_control_inst_n645_51;
wire u_usb_device_controller_n1241_54;
wire u_usb_device_controller_n1242_54;
wire u_usb_device_controller_n1243_54;
wire u_usb_device_controller_n1244_54;
wire u_usb_device_controller_n1241_56;
wire u_usb_device_controller_n1242_56;
wire u_usb_device_controller_n1243_56;
wire u_usb_device_controller_n1244_56;
wire u_usb_device_controller_n1241;
wire u_usb_device_controller_n1242;
wire u_usb_device_controller_n1243;
wire u_usb_device_controller_n1244;
wire u_usb_device_controller_utmi_txvalid_o_d;
wire u_usb_device_controller_n2219;
wire u_usb_device_controller_n384;
wire u_usb_device_controller_n385;
wire u_usb_device_controller_n442;
wire u_usb_device_controller_n443;
wire u_usb_device_controller_n502;
wire u_usb_device_controller_n503;
wire u_usb_device_controller_n560;
wire u_usb_device_controller_n561;
wire u_usb_device_controller_n620;
wire u_usb_device_controller_n621;
wire u_usb_device_controller_n680;
wire u_usb_device_controller_n681;
wire u_usb_device_controller_n742;
wire u_usb_device_controller_n743;
wire u_usb_device_controller_n800;
wire u_usb_device_controller_n801;
wire u_usb_device_controller_n860;
wire u_usb_device_controller_n861;
wire u_usb_device_controller_n920;
wire u_usb_device_controller_n921;
wire u_usb_device_controller_n982;
wire u_usb_device_controller_n983;
wire u_usb_device_controller_n1042;
wire u_usb_device_controller_n1043;
wire u_usb_device_controller_n1104;
wire u_usb_device_controller_n1105;
wire u_usb_device_controller_n1166;
wire u_usb_device_controller_n1167;
wire u_usb_device_controller_n1230;
wire u_usb_device_controller_n1231;
wire u_usb_device_controller_n2339;
wire u_usb_device_controller_txpktfin_o_d;
wire u_usb_device_controller_n2025;
wire u_usb_device_controller_n2026;
wire u_usb_device_controller_n2027;
wire u_usb_device_controller_n2028;
wire u_usb_device_controller_n2029;
wire u_usb_device_controller_n2030;
wire u_usb_device_controller_n2031;
wire u_usb_device_controller_n2032;
wire u_usb_device_controller_n2033;
wire u_usb_device_controller_test_packet_inst_n127;
wire u_usb_device_controller_test_packet_inst_n128;
wire u_usb_device_controller_test_packet_inst_n129;
wire u_usb_device_controller_test_packet_inst_n130;
wire u_usb_device_controller_test_packet_inst_n131;
wire u_usb_device_controller_test_packet_inst_n132;
wire u_usb_device_controller_test_packet_inst_n133;
wire u_usb_device_controller_test_packet_inst_n134;
wire u_usb_device_controller_test_packet_inst_n135;
wire u_usb_device_controller_test_packet_inst_n136;
wire u_usb_device_controller_test_packet_inst_n137;
wire u_usb_device_controller_test_packet_inst_n138;
wire u_usb_device_controller_test_packet_inst_n378;
wire u_usb_device_controller_u_usb_packet_n778;
wire u_usb_device_controller_u_usb_packet_n779;
wire u_usb_device_controller_u_usb_packet_n780;
wire u_usb_device_controller_u_usb_packet_n781;
wire u_usb_device_controller_u_usb_packet_n782;
wire u_usb_device_controller_u_usb_packet_n783;
wire u_usb_device_controller_u_usb_packet_n784;
wire u_usb_device_controller_u_usb_packet_n785;
wire u_usb_device_controller_u_usb_packet_n912;
wire u_usb_device_controller_u_usb_packet_n919;
wire u_usb_device_controller_u_usb_packet_n920;
wire u_usb_device_controller_usb_transact_inst_T_PING;
wire u_usb_device_controller_usb_transact_inst_n1041;
wire u_usb_device_controller_usb_control_inst_n1629;
wire u_usb_device_controller_usb_control_inst_n2896;
wire u_usb_device_controller_u_usb_init_n212;
wire u_usb_device_controller_u_usb_init_n215;
wire u_usb_device_controller_u_usb_init_n216;
wire u_usb_device_controller_usb_control_inst_n435;
wire u_usb_device_controller_usb_control_inst_n436;
wire u_usb_device_controller_usb_control_inst_n437;
wire u_usb_device_controller_usb_control_inst_n438;
wire u_usb_device_controller_usb_control_inst_n439;
wire u_usb_device_controller_usb_control_inst_n440;
wire u_usb_device_controller_usb_control_inst_n441;
wire u_usb_device_controller_usb_control_inst_n442;
wire u_usb_device_controller_u_usb_init_phy_linestate_rst;
wire u_usb_device_controller_u_usb_packet_n328;
wire u_usb_device_controller_usb_control_inst_n1836;
wire u_usb_device_controller_usb_control_inst_n1837;
wire u_usb_device_controller_usb_control_inst_n1864;
wire u_usb_device_controller_usb_control_inst_n2070;
wire u_usb_device_controller_usb_control_inst_n1876;
wire u_usb_device_controller_u_usb_init_n242;
wire u_usb_device_controller_u_usb_init_n280;
wire u_usb_device_controller_u_usb_packet_n800;
wire u_usb_device_controller_rxdat_d0_7;
wire u_usb_device_controller_u_usb_init_s_state_0;
wire u_usb_device_controller_u_usb_packet_crc16_buf_15;
wire u_usb_device_controller_usb_control_inst_s_answerlen_7;
wire u_usb_device_controller_n1619;
wire u_usb_device_controller_u_usb_packet_n615;
wire u_usb_device_controller_u_usb_packet_s_dataout_7;
wire u_usb_device_controller_usb_transact_inst_n1091;
wire u_usb_device_controller_usb_transact_inst_n1074_19;
wire u_usb_device_controller_usb_transact_inst_n1072_15;
wire u_usb_device_controller_usb_transact_inst_n1157_23;
wire u_usb_device_controller_usb_control_inst_n1670;
wire u_usb_device_controller_usb_control_inst_s_answerptr_7_8;
wire u_usb_device_controller_usb_control_inst_s_answerptr_5;
wire u_usb_device_controller_u_usb_packet_s_state_3;
wire u_usb_device_controller_usb_transact_inst_s_sof_11;
wire u_usb_device_controller_usb_transact_inst_s_sendpid_0;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_1;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_2;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_3;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_4;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_5;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_6;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_7;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_8;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_9;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_10;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_11;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_12;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_13;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_14;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_15;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_1;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_2;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_3;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_4;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_5;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_6;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_7;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_8;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_9;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_10;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_11;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_12;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_13;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_14;
wire u_usb_device_controller_usb_control_inst_C_CLROUT_15;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_1;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_2;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_3;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_4;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_5;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_6;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_7;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_8;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_9;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_10;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_11;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_12;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_13;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_14;
wire u_usb_device_controller_usb_control_inst_C_SHLTIN_15;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_1;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_2;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_3;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_4;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_5;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_6;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_7;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_8;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_9;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_10;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_11;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_12;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_13;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_14;
wire u_usb_device_controller_usb_control_inst_C_SHLTOUT_15;
wire u_usb_device_controller_usb_transact_inst_n1068;
wire u_usb_device_controller_u_usb_packet_n640;
wire u_usb_device_controller_u_usb_packet_n642;
wire u_usb_device_controller_u_usb_packet_n644;
wire u_usb_device_controller_u_usb_packet_n646;
wire u_usb_device_controller_u_usb_packet_n650;
wire u_usb_device_controller_u_usb_packet_n652;
wire u_usb_device_controller_usb_transact_inst_n1064;
wire u_usb_device_controller_usb_transact_inst_n1066;
wire u_usb_device_controller_usb_transact_inst_n1074;
wire u_usb_device_controller_usb_transact_inst_n1070;
wire u_usb_device_controller_usb_transact_inst_n1163;
wire u_usb_device_controller_usb_control_inst_n1672;
wire u_usb_device_controller_usb_control_inst_n1678;
wire u_usb_device_controller_usb_control_inst_n1680;
wire u_usb_device_controller_usb_control_inst_n1682;
wire u_usb_device_controller_usb_control_inst_n1684;
wire u_usb_device_controller_usb_control_inst_n1686;
wire u_usb_device_controller_usb_control_inst_n1688;
wire u_usb_device_controller_usb_control_inst_n1690;
wire u_usb_device_controller_usb_control_inst_n1701;
wire u_usb_device_controller_usb_control_inst_n1703;
wire u_usb_device_controller_usb_control_inst_n1705;
wire u_usb_device_controller_usb_control_inst_n1707;
wire u_usb_device_controller_usb_control_inst_n1709;
wire u_usb_device_controller_usb_control_inst_n1711;
wire u_usb_device_controller_usb_control_inst_n1713;
wire u_usb_device_controller_usb_control_inst_n1715;
wire u_usb_device_controller_usb_control_inst_n1717;
wire u_usb_device_controller_usb_control_inst_n1719;
wire u_usb_device_controller_usb_control_inst_n1721;
wire u_usb_device_controller_usb_control_inst_n1723;
wire u_usb_device_controller_usb_control_inst_n1725;
wire u_usb_device_controller_usb_control_inst_n1727;
wire u_usb_device_controller_usb_control_inst_n1729;
wire u_usb_device_controller_usb_control_inst_n1731;
wire u_usb_device_controller_usb_control_inst_n1733;
wire u_usb_device_controller_usb_control_inst_n1735;
wire u_usb_device_controller_usb_control_inst_n1737;
wire u_usb_device_controller_usb_control_inst_n1739;
wire u_usb_device_controller_usb_control_inst_n1741;
wire u_usb_device_controller_usb_control_inst_n1743;
wire u_usb_device_controller_usb_control_inst_n1745;
wire u_usb_device_controller_usb_control_inst_n1747;
wire u_usb_device_controller_usb_control_inst_n1749;
wire u_usb_device_controller_usb_control_inst_n1751;
wire u_usb_device_controller_usb_control_inst_n1753;
wire u_usb_device_controller_usb_control_inst_n1755;
wire u_usb_device_controller_usb_control_inst_n1757;
wire u_usb_device_controller_usb_control_inst_n1759;
wire u_usb_device_controller_usb_control_inst_n1646;
wire u_usb_device_controller_usb_control_inst_n1649;
wire u_usb_device_controller_usb_control_inst_n1652;
wire u_usb_device_controller_usb_control_inst_n1655;
wire u_usb_device_controller_usb_control_inst_n1658;
wire u_usb_device_controller_usb_control_inst_n1661;
wire u_usb_device_controller_usb_control_inst_n1664;
wire u_usb_device_controller_usb_control_inst_n1696;
wire u_usb_device_controller_u_usb_packet_n626;
wire u_usb_device_controller_u_usb_packet_n628;
wire u_usb_device_controller_u_usb_packet_n630;
wire u_usb_device_controller_u_usb_packet_n632;
wire u_usb_device_controller_u_usb_packet_n633;
wire u_usb_device_controller_u_usb_packet_n635;
wire u_usb_device_controller_usb_transact_inst_n1086;
wire u_usb_device_controller_usb_transact_inst_n1088;
wire u_usb_device_controller_usb_transact_inst_n1090;
wire u_usb_device_controller_usb_transact_inst_n1093;
wire u_usb_device_controller_usb_transact_inst_n1095;
wire u_usb_device_controller_usb_transact_inst_n1097;
wire u_usb_device_controller_usb_transact_inst_n1101;
wire u_usb_device_controller_usb_transact_inst_n1103;
wire u_usb_device_controller_usb_transact_inst_n1105;
wire u_usb_device_controller_usb_transact_inst_n1107;
wire u_usb_device_controller_usb_transact_inst_n1109;
wire u_usb_device_controller_usb_transact_inst_n1138;
wire u_usb_device_controller_usb_transact_inst_n1142;
wire u_usb_device_controller_usb_transact_inst_n1144;
wire u_usb_device_controller_usb_transact_inst_n1146;
wire u_usb_device_controller_usb_transact_inst_n1148;
wire u_usb_device_controller_usb_transact_inst_n1150;
wire u_usb_device_controller_usb_transact_inst_n1152;
wire u_usb_device_controller_usb_transact_inst_n1154;
wire u_usb_device_controller_n1615;
wire u_usb_device_controller_usb_transact_inst_n1076;
wire u_usb_device_controller_usb_transact_inst_n1072;
wire u_usb_device_controller_usb_transact_inst_n1157;
wire u_usb_device_controller_usb_transact_inst_n1159;
wire u_usb_device_controller_usb_transact_inst_n1161;
wire u_usb_device_controller_usb_control_inst_n1860;
wire u_usb_device_controller_n1241_60;
wire u_usb_device_controller_n1242_60;
wire u_usb_device_controller_n1243_60;
wire u_usb_device_controller_n1244_60;
wire u_usb_device_controller_n385_6;
wire u_usb_device_controller_n443_6;
wire u_usb_device_controller_n503_6;
wire u_usb_device_controller_n561_6;
wire u_usb_device_controller_n621_6;
wire u_usb_device_controller_n681_6;
wire u_usb_device_controller_n743_6;
wire u_usb_device_controller_n801_6;
wire u_usb_device_controller_n861_6;
wire u_usb_device_controller_n921_6;
wire u_usb_device_controller_n983_6;
wire u_usb_device_controller_n1043_6;
wire u_usb_device_controller_n1105_6;
wire u_usb_device_controller_n1167_6;
wire u_usb_device_controller_n1231_6;
wire u_usb_device_controller_test_packet_inst_cnt_11;
wire u_usb_device_controller_test_packet_inst_test_data_7;
wire u_usb_device_controller_test_packet_inst_test_data_val;
wire u_usb_device_controller_u_usb_init_s_state_1;
wire u_usb_device_controller_u_usb_init_n218;
wire u_usb_device_controller_test_packet_inst_n319;
wire u_usb_device_controller_test_packet_inst_n318;
wire u_usb_device_controller_test_packet_inst_n317;
wire u_usb_device_controller_test_packet_inst_n312;
wire u_usb_device_controller_test_packet_inst_n311;
wire u_usb_device_controller_n1244_62;
wire u_usb_device_controller_n1243_62;
wire u_usb_device_controller_n1242_62;
wire u_usb_device_controller_n1241_62;
wire u_usb_device_controller_u_usb_init_n208;
wire u_usb_device_controller_u_usb_init_n222;
wire u_usb_device_controller_u_usb_init_n221;
wire u_usb_device_controller_u_usb_init_n220;
wire u_usb_device_controller_u_usb_init_n213;
wire u_usb_device_controller_u_usb_init_n219;
wire u_usb_device_controller_n1534;
wire u_usb_device_controller_n1529;
wire u_usb_device_controller_n1524;
wire u_usb_device_controller_n1519;
wire u_usb_device_controller_usbc_dsclen_1;
wire u_usb_device_controller_usbc_dsclen_2;
wire u_usb_device_controller_usbc_dsclen_3;
wire u_usb_device_controller_usbc_dsclen_4;
wire u_usb_device_controller_usbc_dsclen_5;
wire u_usb_device_controller_usbc_dsclen_7;
wire u_usb_device_controller_descrom_start_0;
wire u_usb_device_controller_descrom_start_1;
wire u_usb_device_controller_descrom_start_2;
wire u_usb_device_controller_descrom_start_3;
wire u_usb_device_controller_descrom_start_4;
wire u_usb_device_controller_descrom_start_5;
wire u_usb_device_controller_descrom_start_6;
wire u_usb_device_controller_descrom_start_7;
wire u_usb_device_controller_descrom_start_8;
wire u_usb_device_controller_descrom_start_9;
wire u_usb_device_controller_usb_transact_inst_txpop_o_d;
wire u_usb_device_controller_test_packet_inst_n315;
wire u_usb_device_controller_test_packet_inst_n313;
wire u_usb_device_controller_test_packet_inst_n316;
wire u_usb_device_controller_test_packet_inst_n314;
wire u_usb_device_controller_u_usb_init_n211;
wire u_usb_device_controller_usb_control_inst_n414;
wire u_usb_device_controller_usb_control_inst_n413;
wire u_usb_device_controller_usb_control_inst_n412;
wire u_usb_device_controller_usb_control_inst_n411;
wire u_usb_device_controller_usb_control_inst_n410;
wire u_usb_device_controller_usb_control_inst_n409;
wire u_usb_device_controller_usb_control_inst_n408;
wire u_usb_device_controller_usb_control_inst_n407;
wire u_usb_device_controller_u_usb_packet_n776;
wire u_usb_device_controller_u_usb_packet_n775;
wire u_usb_device_controller_u_usb_packet_n764;
wire u_usb_device_controller_u_usb_packet_n761;
wire u_usb_device_controller_u_usb_init_n217;
wire u_usb_device_controller_n1261;
wire u_usb_device_controller_u_usb_packet_crc5_buf_4;
wire u_usb_device_controller_usb_control_inst_s_answerptr_7;
wire u_usb_device_controller_usb_control_inst_s_sendbyte_1;
wire u_usb_device_controller_s_nyet_9;
wire u_usb_device_controller_usb_transact_inst_s_sof_valid;
wire u_usb_device_controller_n1581;
wire u_usb_device_controller_usb_control_inst_n1388;
wire u_usb_device_controller_usb_control_inst_n1387;
wire u_usb_device_controller_usb_control_inst_n1386;
wire u_usb_device_controller_usb_control_inst_n1385;
wire u_usb_device_controller_usb_control_inst_n1384;
wire u_usb_device_controller_usb_control_inst_n1383;
wire u_usb_device_controller_usb_control_inst_n1382;
wire u_usb_device_controller_usb_control_inst_n1617;
wire u_usb_device_controller_usb_transact_inst_n1136;
wire u_usb_device_controller_usb_transact_inst_n1133;
wire u_usb_device_controller_usb_transact_inst_n1130;
wire u_usb_device_controller_usb_transact_inst_n1127;
wire u_usb_device_controller_usb_transact_inst_n1124;
wire u_usb_device_controller_usb_transact_inst_n1121;
wire u_usb_device_controller_usb_transact_inst_n1118;
wire u_usb_device_controller_n1609;
wire u_usb_device_controller_n1605;
wire u_usb_device_controller_n1603;
wire u_usb_device_controller_n1599;
wire u_usb_device_controller_n1597;
wire u_usb_device_controller_n1593;
wire u_usb_device_controller_u_usb_packet_n579;
wire u_usb_device_controller_u_usb_packet_n577;
wire u_usb_device_controller_u_usb_packet_n575;
wire u_usb_device_controller_u_usb_packet_n573;
wire u_usb_device_controller_u_usb_packet_n571;
wire u_usb_device_controller_utmi_dataout_o_d_7;
wire u_usb_device_controller_utmi_dataout_o_d_6;
wire u_usb_device_controller_utmi_dataout_o_d_5;
wire u_usb_device_controller_utmi_dataout_o_d_4;
wire u_usb_device_controller_utmi_dataout_o_d_3;
wire u_usb_device_controller_utmi_dataout_o_d_2;
wire u_usb_device_controller_utmi_dataout_o_d_1;
wire u_usb_device_controller_utmi_dataout_o_d_0;
wire u_usb_device_controller_rxact_o_d_3;
wire u_usb_device_controller_n2339_4;
wire u_usb_device_controller_n1585_4;
wire u_usb_device_controller_setup_o_d_3;
wire u_usb_device_controller_n2024_4;
wire u_usb_device_controller_test_packet_inst_n127_6;
wire u_usb_device_controller_test_packet_inst_n127_7;
wire u_usb_device_controller_test_packet_inst_n129_6;
wire u_usb_device_controller_test_packet_inst_n130_6;
wire u_usb_device_controller_test_packet_inst_n133_6;
wire u_usb_device_controller_test_packet_inst_n133_7;
wire u_usb_device_controller_test_packet_inst_n378_4;
wire u_usb_device_controller_u_usb_init_n414_4;
wire u_usb_device_controller_u_usb_packet_n782_4;
wire u_usb_device_controller_u_usb_packet_n782_5;
wire u_usb_device_controller_u_usb_packet_n784_4;
wire u_usb_device_controller_u_usb_packet_n784_6;
wire u_usb_device_controller_u_usb_packet_n785_4;
wire u_usb_device_controller_u_usb_packet_n785_5;
wire u_usb_device_controller_u_usb_packet_n912_4;
wire u_usb_device_controller_u_usb_packet_n912_5;
wire u_usb_device_controller_u_usb_packet_n912_6;
wire u_usb_device_controller_u_usb_packet_n912_7;
wire u_usb_device_controller_u_usb_packet_n920_4;
wire u_usb_device_controller_usb_transact_inst_n1041_4;
wire u_usb_device_controller_usb_transact_inst_n1041_6;
wire u_usb_device_controller_usb_transact_inst_n1565_4;
wire u_usb_device_controller_usb_transact_inst_n1565_5;
wire u_usb_device_controller_usb_control_inst_n1629_4;
wire u_usb_device_controller_usb_control_inst_n1629_5;
wire u_usb_device_controller_usb_control_inst_n1629_6;
wire u_usb_device_controller_usb_control_inst_n2896_4;
wire u_usb_device_controller_usb_control_inst_n2896_5;
wire u_usb_device_controller_u_usb_init_n212_28;
wire u_usb_device_controller_u_usb_init_n212_29;
wire u_usb_device_controller_u_usb_init_n212_31;
wire u_usb_device_controller_u_usb_init_n215_52;
wire u_usb_device_controller_u_usb_init_n216_49;
wire u_usb_device_controller_u_usb_init_n216_51;
wire u_usb_device_controller_usb_control_inst_n435_16;
wire u_usb_device_controller_usb_control_inst_n435_17;
wire u_usb_device_controller_u_usb_packet_n328_10;
wire u_usb_device_controller_u_usb_packet_n328_11;
wire u_usb_device_controller_usb_control_inst_n1836_8;
wire u_usb_device_controller_usb_control_inst_n1837_6;
wire u_usb_device_controller_usb_control_inst_n1837_7;
wire u_usb_device_controller_usb_control_inst_n2067_6;
wire u_usb_device_controller_usb_control_inst_n2067_7;
wire u_usb_device_controller_u_usb_packet_n800_6;
wire u_usb_device_controller_rxdat_d0_7_9;
wire u_usb_device_controller_rxdat_d0_7_10;
wire u_usb_device_controller_u_usb_init_s_opmode_1;
wire u_usb_device_controller_u_usb_init_s_state_3;
wire u_usb_device_controller_u_usb_init_s_state_3_10;
wire u_usb_device_controller_u_usb_init_s_chirpcnt_2_8;
wire u_usb_device_controller_usb_control_inst_s_answerlen_7_7;
wire u_usb_device_controller_u_usb_packet_n615_42;
wire u_usb_device_controller_u_usb_packet_s_dataout_7_9;
wire u_usb_device_controller_usb_transact_inst_n1080;
wire u_usb_device_controller_usb_transact_inst_n1080_46;
wire u_usb_device_controller_usb_transact_inst_n1064_16;
wire u_usb_device_controller_usb_transact_inst_n1074_22;
wire u_usb_device_controller_usb_transact_inst_n1072_18;
wire u_usb_device_controller_usb_transact_inst_n1072_19;
wire u_usb_device_controller_usb_transact_inst_n1138_24;
wire u_usb_device_controller_usb_transact_inst_n1138_25;
wire u_usb_device_controller_usb_transact_inst_n1157_26;
wire u_usb_device_controller_usb_transact_inst_n1157_27;
wire u_usb_device_controller_usb_transact_inst_n1157_28;
wire u_usb_device_controller_usb_transact_inst_n1157_29;
wire u_usb_device_controller_usb_control_inst_n1670_39;
wire u_usb_device_controller_usb_control_inst_n1670_40;
wire u_usb_device_controller_usb_control_inst_n1670_41;
wire u_usb_device_controller_usb_control_inst_s_answerptr_7_11;
wire u_usb_device_controller_usb_control_inst_s_answerptr_7_12;
wire u_usb_device_controller_usb_control_inst_s_answerptr_5_10;
wire u_usb_device_controller_usb_control_inst_s_sendbyte_7_13;
wire u_usb_device_controller_u_usb_packet_s_state_11;
wire u_usb_device_controller_usb_transact_inst_s_sendpid_3_11;
wire u_usb_device_controller_usb_transact_inst_n1068_10;
wire u_usb_device_controller_u_usb_packet_n640_18;
wire u_usb_device_controller_u_usb_packet_n640_19;
wire u_usb_device_controller_u_usb_packet_n642_18;
wire u_usb_device_controller_u_usb_packet_n642_19;
wire u_usb_device_controller_u_usb_packet_n642_20;
wire u_usb_device_controller_u_usb_packet_n644_18;
wire u_usb_device_controller_u_usb_packet_n644_19;
wire u_usb_device_controller_u_usb_packet_n644_20;
wire u_usb_device_controller_u_usb_packet_n646_18;
wire u_usb_device_controller_u_usb_packet_n646_19;
wire u_usb_device_controller_u_usb_packet_n650_18;
wire u_usb_device_controller_u_usb_packet_n650_19;
wire u_usb_device_controller_u_usb_packet_n652_18;
wire u_usb_device_controller_u_usb_packet_n654_18;
wire u_usb_device_controller_usb_transact_inst_n1064_18;
wire u_usb_device_controller_usb_transact_inst_n1066_14;
wire u_usb_device_controller_usb_transact_inst_n1111_18;
wire u_usb_device_controller_usb_transact_inst_n1074_23;
wire u_usb_device_controller_usb_transact_inst_n1074_24;
wire u_usb_device_controller_usb_transact_inst_n1070_14;
wire u_usb_device_controller_usb_control_inst_n1672_41;
wire u_usb_device_controller_usb_control_inst_n1672_42;
wire u_usb_device_controller_usb_control_inst_n1672_43;
wire u_usb_device_controller_usb_control_inst_n1672_44;
wire u_usb_device_controller_usb_control_inst_n1674_39;
wire u_usb_device_controller_usb_control_inst_n1676_39;
wire u_usb_device_controller_usb_control_inst_n1678_40;
wire u_usb_device_controller_usb_control_inst_n1678_41;
wire u_usb_device_controller_usb_control_inst_n1680_42;
wire u_usb_device_controller_usb_control_inst_n1680_43;
wire u_usb_device_controller_usb_control_inst_n1680_44;
wire u_usb_device_controller_usb_control_inst_n1682_39;
wire u_usb_device_controller_usb_control_inst_n1682_40;
wire u_usb_device_controller_usb_control_inst_n1684_39;
wire u_usb_device_controller_usb_control_inst_n1684_40;
wire u_usb_device_controller_usb_control_inst_n1686_39;
wire u_usb_device_controller_usb_control_inst_n1686_40;
wire u_usb_device_controller_usb_control_inst_n1688_39;
wire u_usb_device_controller_usb_control_inst_n1690_34;
wire u_usb_device_controller_usb_control_inst_n1690_35;
wire u_usb_device_controller_usb_control_inst_n1690_36;
wire u_usb_device_controller_usb_control_inst_n1701_16;
wire u_usb_device_controller_usb_control_inst_n1701_17;
wire u_usb_device_controller_usb_control_inst_n1701_18;
wire u_usb_device_controller_usb_control_inst_n1703_16;
wire u_usb_device_controller_usb_control_inst_n1705_16;
wire u_usb_device_controller_usb_control_inst_n1707_16;
wire u_usb_device_controller_usb_control_inst_n1711_16;
wire u_usb_device_controller_usb_control_inst_n1713_16;
wire u_usb_device_controller_usb_control_inst_n1715_16;
wire u_usb_device_controller_usb_control_inst_n1715_17;
wire u_usb_device_controller_usb_control_inst_n1731_16;
wire u_usb_device_controller_usb_control_inst_n1745_16;
wire u_usb_device_controller_usb_control_inst_n1775_13;
wire u_usb_device_controller_usb_control_inst_n1805_13;
wire u_usb_device_controller_usb_control_inst_n1649_16;
wire u_usb_device_controller_usb_control_inst_n1649_17;
wire u_usb_device_controller_usb_control_inst_n1649_18;
wire u_usb_device_controller_usb_control_inst_n1652_16;
wire u_usb_device_controller_usb_control_inst_n1652_18;
wire u_usb_device_controller_usb_control_inst_n1658_16;
wire u_usb_device_controller_usb_control_inst_n1661_16;
wire u_usb_device_controller_usb_control_inst_n1661_17;
wire u_usb_device_controller_usb_control_inst_n1661_18;
wire u_usb_device_controller_usb_control_inst_n1661_19;
wire u_usb_device_controller_u_usb_packet_n620_47;
wire u_usb_device_controller_u_usb_packet_n626_41;
wire u_usb_device_controller_u_usb_packet_n626_42;
wire u_usb_device_controller_u_usb_packet_n628_47;
wire u_usb_device_controller_u_usb_packet_n633_39;
wire u_usb_device_controller_usb_transact_inst_n1088_44;
wire u_usb_device_controller_usb_transact_inst_n1088_45;
wire u_usb_device_controller_usb_transact_inst_n1090_46;
wire u_usb_device_controller_usb_transact_inst_n1091_49;
wire u_usb_device_controller_usb_transact_inst_n1091_50;
wire u_usb_device_controller_usb_transact_inst_n1093_51;
wire u_usb_device_controller_usb_transact_inst_n1095_44;
wire u_usb_device_controller_usb_transact_inst_n1095_45;
wire u_usb_device_controller_usb_transact_inst_n1095_46;
wire u_usb_device_controller_usb_transact_inst_n1099_47;
wire u_usb_device_controller_usb_transact_inst_n1101_44;
wire u_usb_device_controller_usb_transact_inst_n1105_47;
wire u_usb_device_controller_usb_transact_inst_n1105_48;
wire u_usb_device_controller_usb_transact_inst_n1109_47;
wire u_usb_device_controller_usb_transact_inst_n1109_48;
wire u_usb_device_controller_usb_transact_inst_n1138_29;
wire u_usb_device_controller_usb_transact_inst_n1138_30;
wire u_usb_device_controller_usb_transact_inst_n1140_22;
wire u_usb_device_controller_usb_transact_inst_n1142_23;
wire u_usb_device_controller_usb_transact_inst_n1144_22;
wire u_usb_device_controller_usb_transact_inst_n1146_22;
wire u_usb_device_controller_usb_transact_inst_n1148_22;
wire u_usb_device_controller_usb_transact_inst_n1150_22;
wire u_usb_device_controller_usb_transact_inst_n1152_22;
wire u_usb_device_controller_n1615_15;
wire u_usb_device_controller_usb_transact_inst_n1076_21;
wire u_usb_device_controller_usb_transact_inst_n1072_20;
wire u_usb_device_controller_usb_transact_inst_n1157_30;
wire u_usb_device_controller_usb_transact_inst_n1157_31;
wire u_usb_device_controller_usb_transact_inst_n1159_25;
wire u_usb_device_controller_usb_transact_inst_n1159_26;
wire u_usb_device_controller_usb_control_inst_n1860_29;
wire u_usb_device_controller_usb_control_inst_n1860_30;
wire u_usb_device_controller_n385_7;
wire u_usb_device_controller_n443_7;
wire u_usb_device_controller_n503_7;
wire u_usb_device_controller_n561_7;
wire u_usb_device_controller_usb_control_inst_s_ctlparam_7_7;
wire u_usb_device_controller_isync_1_10;
wire u_usb_device_controller_isync_2_9;
wire u_usb_device_controller_isync_3_9;
wire u_usb_device_controller_isync_4_10;
wire u_usb_device_controller_test_packet_inst_cnt_11_9;
wire u_usb_device_controller_test_packet_inst_cnt_11_10;
wire u_usb_device_controller_test_packet_inst_test_data_6;
wire u_usb_device_controller_test_packet_inst_test_data_6_8;
wire u_usb_device_controller_u_usb_init_s_state_2_14;
wire u_usb_device_controller_test_packet_inst_n318_8;
wire u_usb_device_controller_test_packet_inst_n318_9;
wire u_usb_device_controller_test_packet_inst_n318_10;
wire u_usb_device_controller_test_packet_inst_n317_9;
wire u_usb_device_controller_test_packet_inst_n317_10;
wire u_usb_device_controller_test_packet_inst_n312_8;
wire u_usb_device_controller_test_packet_inst_n312_9;
wire u_usb_device_controller_test_packet_inst_n312_10;
wire u_usb_device_controller_test_packet_inst_n311_9;
wire u_usb_device_controller_u_usb_init_n213_28;
wire u_usb_device_controller_u_usb_init_n219_28;
wire u_usb_device_controller_n1534_26;
wire u_usb_device_controller_n1534_28;
wire u_usb_device_controller_n1534_29;
wire u_usb_device_controller_n1529_24;
wire u_usb_device_controller_n1529_25;
wire u_usb_device_controller_n1529_26;
wire u_usb_device_controller_n1524_25;
wire u_usb_device_controller_usbc_dsclen_0_15;
wire u_usb_device_controller_usbc_dsclen_1_14;
wire u_usb_device_controller_usbc_dsclen_1_15;
wire u_usb_device_controller_usbc_dsclen_2_14;
wire u_usb_device_controller_usbc_dsclen_2_15;
wire u_usb_device_controller_usbc_dsclen_3_14;
wire u_usb_device_controller_usbc_dsclen_4_14;
wire u_usb_device_controller_usbc_dsclen_4_15;
wire u_usb_device_controller_usbc_dsclen_5_14;
wire u_usb_device_controller_usbc_dsclen_6_14;
wire u_usb_device_controller_usbc_dsclen_6_15;
wire u_usb_device_controller_usbc_dsclen_7_14;
wire u_usb_device_controller_descrom_start_0_14;
wire u_usb_device_controller_descrom_start_0_15;
wire u_usb_device_controller_descrom_start_1_14;
wire u_usb_device_controller_descrom_start_1_15;
wire u_usb_device_controller_descrom_start_2_14;
wire u_usb_device_controller_descrom_start_2_15;
wire u_usb_device_controller_descrom_start_3_14;
wire u_usb_device_controller_descrom_start_3_15;
wire u_usb_device_controller_descrom_start_4_14;
wire u_usb_device_controller_descrom_start_4_15;
wire u_usb_device_controller_descrom_start_5_14;
wire u_usb_device_controller_descrom_start_5_15;
wire u_usb_device_controller_descrom_start_6_14;
wire u_usb_device_controller_descrom_start_6_15;
wire u_usb_device_controller_descrom_start_7_14;
wire u_usb_device_controller_descrom_start_7_15;
wire u_usb_device_controller_descrom_start_8_14;
wire u_usb_device_controller_descrom_start_8_15;
wire u_usb_device_controller_descrom_start_9_14;
wire u_usb_device_controller_descrom_start_9_15;
wire u_usb_device_controller_usb_transact_inst_txpop_o_d_5;
wire u_usb_device_controller_test_packet_inst_n313_8;
wire u_usb_device_controller_test_packet_inst_n316_8;
wire u_usb_device_controller_test_packet_inst_n314_8;
wire u_usb_device_controller_test_packet_inst_n314_9;
wire u_usb_device_controller_n1810_6;
wire u_usb_device_controller_u_usb_packet_n776_6;
wire u_usb_device_controller_u_usb_packet_n776_7;
wire u_usb_device_controller_u_usb_packet_n776_8;
wire u_usb_device_controller_u_usb_packet_n776_9;
wire u_usb_device_controller_u_usb_packet_n775_6;
wire u_usb_device_controller_u_usb_packet_n775_7;
wire u_usb_device_controller_u_usb_packet_n775_8;
wire u_usb_device_controller_u_usb_packet_n774_6;
wire u_usb_device_controller_u_usb_packet_n774_7;
wire u_usb_device_controller_u_usb_packet_n771_6;
wire u_usb_device_controller_u_usb_packet_n771_7;
wire u_usb_device_controller_u_usb_packet_n770_6;
wire u_usb_device_controller_u_usb_packet_n767_6;
wire u_usb_device_controller_u_usb_packet_n761_6;
wire u_usb_device_controller_u_usb_init_n217_37;
wire u_usb_device_controller_u_usb_init_n217_38;
wire u_usb_device_controller_usb_control_inst_usbc_dscrd_4;
wire u_usb_device_controller_usb_control_inst_s_answerptr_7_13;
wire u_usb_device_controller_usb_control_inst_s_sendbyte_7_14;
wire u_usb_device_controller_usb_control_inst_s_interface_set_8;
wire u_usb_device_controller_usb_control_inst_s_interface_set_9;
wire u_usb_device_controller_usb_transact_inst_n1133_26;
wire u_usb_device_controller_usb_transact_inst_n1127_26;
wire u_usb_device_controller_usb_transact_inst_n1118_26;
wire u_usb_device_controller_n1613_21;
wire u_usb_device_controller_n1611_21;
wire u_usb_device_controller_n1603_21;
wire u_usb_device_controller_n1597_21;
wire u_usb_device_controller_u_usb_packet_n579_19;
wire u_usb_device_controller_u_usb_packet_n579_20;
wire u_usb_device_controller_u_usb_packet_n577_19;
wire u_usb_device_controller_u_usb_packet_n577_20;
wire u_usb_device_controller_u_usb_packet_n575_19;
wire u_usb_device_controller_u_usb_packet_n573_19;
wire u_usb_device_controller_u_usb_packet_n571_19;
wire u_usb_device_controller_utmi_dataout_o_d_7_7;
wire u_usb_device_controller_utmi_dataout_o_d_0_4;
wire u_usb_device_controller_utmi_dataout_o_d_0_5;
wire u_usb_device_controller_n2339_5;
wire u_usb_device_controller_n2339_6;
wire u_usb_device_controller_n2024_5;
wire u_usb_device_controller_n2024_6;
wire u_usb_device_controller_test_packet_inst_n130_7;
wire u_usb_device_controller_test_packet_inst_n378_5;
wire u_usb_device_controller_u_usb_packet_n782_6;
wire u_usb_device_controller_u_usb_packet_n782_7;
wire u_usb_device_controller_u_usb_packet_n782_8;
wire u_usb_device_controller_u_usb_packet_n782_9;
wire u_usb_device_controller_u_usb_packet_n784_7;
wire u_usb_device_controller_u_usb_packet_n784_8;
wire u_usb_device_controller_u_usb_packet_n784_9;
wire u_usb_device_controller_u_usb_packet_n784_10;
wire u_usb_device_controller_u_usb_packet_n784_11;
wire u_usb_device_controller_u_usb_packet_n785_6;
wire u_usb_device_controller_u_usb_packet_n785_7;
wire u_usb_device_controller_u_usb_packet_n1454_5;
wire u_usb_device_controller_u_usb_packet_n912_8;
wire u_usb_device_controller_u_usb_packet_n912_9;
wire u_usb_device_controller_u_usb_packet_n912_10;
wire u_usb_device_controller_u_usb_packet_n912_11;
wire u_usb_device_controller_u_usb_packet_n912_12;
wire u_usb_device_controller_u_usb_packet_n912_13;
wire u_usb_device_controller_u_usb_packet_n919_5;
wire u_usb_device_controller_u_usb_packet_n920_6;
wire u_usb_device_controller_u_usb_packet_n920_7;
wire u_usb_device_controller_usb_transact_inst_n1565_7;
wire u_usb_device_controller_usb_control_inst_n2902_5;
wire u_usb_device_controller_u_usb_init_n212_33;
wire u_usb_device_controller_u_usb_init_n212_35;
wire u_usb_device_controller_u_usb_init_n212_37;
wire u_usb_device_controller_u_usb_init_n212_38;
wire u_usb_device_controller_u_usb_init_n212_39;
wire u_usb_device_controller_u_usb_init_n215_53;
wire u_usb_device_controller_u_usb_init_n215_54;
wire u_usb_device_controller_u_usb_init_n215_57;
wire u_usb_device_controller_u_usb_init_n216_52;
wire u_usb_device_controller_u_usb_init_n216_53;
wire u_usb_device_controller_u_usb_init_n216_54;
wire u_usb_device_controller_usb_control_inst_n435_18;
wire u_usb_device_controller_usb_control_inst_n435_19;
wire u_usb_device_controller_usb_control_inst_n435_20;
wire u_usb_device_controller_u_usb_packet_n328_12;
wire u_usb_device_controller_u_usb_packet_n328_13;
wire u_usb_device_controller_u_usb_packet_n328_14;
wire u_usb_device_controller_u_usb_packet_n328_16;
wire u_usb_device_controller_u_usb_packet_n328_17;
wire u_usb_device_controller_usb_control_inst_n1836_9;
wire u_usb_device_controller_usb_control_inst_n1836_10;
wire u_usb_device_controller_usb_transact_inst_s_endpt_0_7;
wire u_usb_device_controller_u_usb_init_s_state_3_11;
wire u_usb_device_controller_u_usb_init_s_state_3_12;
wire u_usb_device_controller_u_usb_init_s_chirpcnt_2_9;
wire u_usb_device_controller_u_usb_init_s_chirpcnt_2_10;
wire u_usb_device_controller_u_usb_packet_n615_43;
wire u_usb_device_controller_u_usb_packet_n615_44;
wire u_usb_device_controller_u_usb_packet_n615_45;
wire u_usb_device_controller_u_usb_packet_n615_46;
wire u_usb_device_controller_usb_transact_inst_n1080_48;
wire u_usb_device_controller_usb_transact_inst_n1080_49;
wire u_usb_device_controller_usb_transact_inst_n1064_20;
wire u_usb_device_controller_usb_transact_inst_n1074_25;
wire u_usb_device_controller_usb_transact_inst_n1072_21;
wire u_usb_device_controller_usb_control_inst_n1670_43;
wire u_usb_device_controller_usb_control_inst_s_answerptr_7_14;
wire u_usb_device_controller_usb_control_inst_s_answerptr_7_15;
wire u_usb_device_controller_usb_control_inst_s_answerptr_5_12;
wire u_usb_device_controller_usb_control_inst_s_sendbyte_7_15;
wire u_usb_device_controller_usb_control_inst_s_sendbyte_7_16;
wire u_usb_device_controller_u_usb_packet_s_state_11_21;
wire u_usb_device_controller_u_usb_packet_s_state_11_22;
wire u_usb_device_controller_u_usb_packet_s_state_11_23;
wire u_usb_device_controller_usb_transact_inst_s_sendpid_3_13;
wire u_usb_device_controller_usb_transact_inst_s_sendpid_3_14;
wire u_usb_device_controller_u_usb_packet_n640_21;
wire u_usb_device_controller_u_usb_packet_n642_21;
wire u_usb_device_controller_u_usb_packet_n644_21;
wire u_usb_device_controller_u_usb_packet_n646_20;
wire u_usb_device_controller_u_usb_packet_n650_20;
wire u_usb_device_controller_u_usb_packet_n650_21;
wire u_usb_device_controller_usb_transact_inst_n1064_21;
wire u_usb_device_controller_usb_control_inst_n1672_45;
wire u_usb_device_controller_usb_control_inst_n1672_46;
wire u_usb_device_controller_usb_control_inst_n1678_42;
wire u_usb_device_controller_usb_control_inst_n1678_43;
wire u_usb_device_controller_usb_control_inst_n1678_44;
wire u_usb_device_controller_usb_control_inst_n1680_46;
wire u_usb_device_controller_usb_control_inst_n1680_47;
wire u_usb_device_controller_usb_control_inst_n1684_41;
wire u_usb_device_controller_usb_control_inst_n1684_42;
wire u_usb_device_controller_usb_control_inst_n1686_41;
wire u_usb_device_controller_usb_control_inst_n1686_42;
wire u_usb_device_controller_usb_control_inst_n1690_37;
wire u_usb_device_controller_usb_control_inst_n1690_38;
wire u_usb_device_controller_usb_control_inst_n1709_17;
wire u_usb_device_controller_usb_control_inst_n1649_19;
wire u_usb_device_controller_usb_control_inst_n1649_21;
wire u_usb_device_controller_usb_control_inst_n1652_19;
wire u_usb_device_controller_u_usb_packet_n626_44;
wire u_usb_device_controller_u_usb_packet_n626_45;
wire u_usb_device_controller_u_usb_packet_n626_46;
wire u_usb_device_controller_u_usb_packet_n628_48;
wire u_usb_device_controller_u_usb_packet_n633_40;
wire u_usb_device_controller_u_usb_packet_n633_41;
wire u_usb_device_controller_u_usb_packet_n633_42;
wire u_usb_device_controller_usb_transact_inst_n1091_52;
wire u_usb_device_controller_usb_transact_inst_n1095_47;
wire u_usb_device_controller_usb_transact_inst_n1101_45;
wire u_usb_device_controller_usb_transact_inst_n1109_49;
wire u_usb_device_controller_usb_transact_inst_n1138_31;
wire u_usb_device_controller_usb_transact_inst_n1072_22;
wire u_usb_device_controller_usb_transact_inst_n1159_27;
wire u_usb_device_controller_usb_control_inst_n1860_31;
wire u_usb_device_controller_usb_control_inst_n1860_32;
wire u_usb_device_controller_usb_control_inst_s_ctlparam_7_8;
wire u_usb_device_controller_test_packet_inst_cnt_11_11;
wire u_usb_device_controller_test_packet_inst_cnt_11_12;
wire u_usb_device_controller_test_packet_inst_cnt_11_13;
wire u_usb_device_controller_test_packet_inst_test_data_6_9;
wire u_usb_device_controller_u_usb_init_s_state_2_16;
wire u_usb_device_controller_test_packet_inst_n318_11;
wire u_usb_device_controller_test_packet_inst_n318_12;
wire u_usb_device_controller_test_packet_inst_n318_13;
wire u_usb_device_controller_test_packet_inst_n318_14;
wire u_usb_device_controller_test_packet_inst_n317_11;
wire u_usb_device_controller_test_packet_inst_n311_10;
wire u_usb_device_controller_u_usb_init_n219_29;
wire u_usb_device_controller_n1534_30;
wire u_usb_device_controller_n1534_31;
wire u_usb_device_controller_n1534_32;
wire u_usb_device_controller_n1534_33;
wire u_usb_device_controller_n1534_34;
wire u_usb_device_controller_n1529_28;
wire u_usb_device_controller_n1529_29;
wire u_usb_device_controller_usbc_dsclen_0_16;
wire u_usb_device_controller_usbc_dsclen_0_17;
wire u_usb_device_controller_usbc_dsclen_0_18;
wire u_usb_device_controller_usbc_dsclen_0_19;
wire u_usb_device_controller_usbc_dsclen_1_16;
wire u_usb_device_controller_usbc_dsclen_1_18;
wire u_usb_device_controller_usbc_dsclen_1_20;
wire u_usb_device_controller_usbc_dsclen_2_16;
wire u_usb_device_controller_usbc_dsclen_2_17;
wire u_usb_device_controller_usbc_dsclen_3_15;
wire u_usb_device_controller_usbc_dsclen_3_16;
wire u_usb_device_controller_usbc_dsclen_3_17;
wire u_usb_device_controller_usbc_dsclen_4_16;
wire u_usb_device_controller_usbc_dsclen_4_17;
wire u_usb_device_controller_usbc_dsclen_4_18;
wire u_usb_device_controller_usbc_dsclen_5_15;
wire u_usb_device_controller_usbc_dsclen_5_16;
wire u_usb_device_controller_usbc_dsclen_5_17;
wire u_usb_device_controller_usbc_dsclen_6_16;
wire u_usb_device_controller_usbc_dsclen_6_17;
wire u_usb_device_controller_usbc_dsclen_7_15;
wire u_usb_device_controller_usbc_dsclen_7_16;
wire u_usb_device_controller_usbc_dsclen_7_17;
wire u_usb_device_controller_descrom_start_0_16;
wire u_usb_device_controller_descrom_start_0_17;
wire u_usb_device_controller_descrom_start_0_18;
wire u_usb_device_controller_descrom_start_1_16;
wire u_usb_device_controller_descrom_start_1_17;
wire u_usb_device_controller_descrom_start_1_18;
wire u_usb_device_controller_descrom_start_2_16;
wire u_usb_device_controller_descrom_start_2_17;
wire u_usb_device_controller_descrom_start_2_18;
wire u_usb_device_controller_descrom_start_3_16;
wire u_usb_device_controller_descrom_start_3_17;
wire u_usb_device_controller_descrom_start_3_18;
wire u_usb_device_controller_descrom_start_4_16;
wire u_usb_device_controller_descrom_start_4_17;
wire u_usb_device_controller_descrom_start_4_18;
wire u_usb_device_controller_descrom_start_5_16;
wire u_usb_device_controller_descrom_start_5_17;
wire u_usb_device_controller_descrom_start_5_18;
wire u_usb_device_controller_descrom_start_6_16;
wire u_usb_device_controller_descrom_start_6_17;
wire u_usb_device_controller_descrom_start_6_18;
wire u_usb_device_controller_descrom_start_7_16;
wire u_usb_device_controller_descrom_start_7_17;
wire u_usb_device_controller_descrom_start_7_18;
wire u_usb_device_controller_descrom_start_8_16;
wire u_usb_device_controller_descrom_start_8_17;
wire u_usb_device_controller_descrom_start_8_18;
wire u_usb_device_controller_descrom_start_9_16;
wire u_usb_device_controller_descrom_start_9_17;
wire u_usb_device_controller_descrom_start_9_18;
wire u_usb_device_controller_usb_transact_inst_txpop_o_d_7;
wire u_usb_device_controller_test_packet_inst_n313_9;
wire u_usb_device_controller_u_usb_packet_n774_8;
wire u_usb_device_controller_u_usb_packet_n774_9;
wire u_usb_device_controller_u_usb_packet_n774_10;
wire u_usb_device_controller_u_usb_packet_n774_11;
wire u_usb_device_controller_u_usb_packet_n771_8;
wire u_usb_device_controller_u_usb_packet_n771_9;
wire u_usb_device_controller_u_usb_packet_n771_10;
wire u_usb_device_controller_u_usb_packet_n771_11;
wire u_usb_device_controller_u_usb_packet_n771_12;
wire u_usb_device_controller_u_usb_packet_n767_8;
wire u_usb_device_controller_u_usb_packet_crc5_buf_4_11;
wire u_usb_device_controller_usb_transact_inst_n1133_27;
wire u_usb_device_controller_u_usb_packet_n579_21;
wire u_usb_device_controller_u_usb_packet_n579_22;
wire u_usb_device_controller_utmi_dataout_o_d_7_8;
wire u_usb_device_controller_n2024_7;
wire u_usb_device_controller_u_usb_packet_n784_13;
wire u_usb_device_controller_u_usb_packet_n785_8;
wire u_usb_device_controller_u_usb_packet_n912_14;
wire u_usb_device_controller_u_usb_packet_n912_15;
wire u_usb_device_controller_u_usb_packet_n912_16;
wire u_usb_device_controller_u_usb_packet_n912_17;
wire u_usb_device_controller_u_usb_packet_n912_18;
wire u_usb_device_controller_u_usb_packet_n912_19;
wire u_usb_device_controller_u_usb_packet_n912_20;
wire u_usb_device_controller_u_usb_packet_n912_21;
wire u_usb_device_controller_usb_control_inst_n2896_7;
wire u_usb_device_controller_u_usb_init_n212_41;
wire u_usb_device_controller_u_usb_init_n212_42;
wire u_usb_device_controller_u_usb_init_n212_43;
wire u_usb_device_controller_u_usb_init_n212_44;
wire u_usb_device_controller_u_usb_init_n212_45;
wire u_usb_device_controller_u_usb_init_n215_58;
wire u_usb_device_controller_u_usb_init_n215_59;
wire u_usb_device_controller_u_usb_packet_n328_20;
wire u_usb_device_controller_u_usb_packet_n328_21;
wire u_usb_device_controller_u_usb_packet_n328_22;
wire u_usb_device_controller_u_usb_packet_n328_23;
wire u_usb_device_controller_u_usb_packet_n328_24;
wire u_usb_device_controller_usb_control_inst_n1836_11;
wire u_usb_device_controller_u_usb_init_s_state_3_13;
wire u_usb_device_controller_u_usb_init_s_state_3_14;
wire u_usb_device_controller_u_usb_init_s_chirpcnt_2_11;
wire u_usb_device_controller_u_usb_init_s_chirpcnt_2_12;
wire u_usb_device_controller_u_usb_init_s_chirpcnt_2_13;
wire u_usb_device_controller_u_usb_init_s_chirpcnt_2_14;
wire u_usb_device_controller_u_usb_packet_n615_47;
wire u_usb_device_controller_usb_control_inst_s_answerptr_7_16;
wire u_usb_device_controller_usb_control_inst_s_sendbyte_7_17;
wire u_usb_device_controller_u_usb_packet_s_state_11_25;
wire u_usb_device_controller_usb_transact_inst_s_sendpid_3_16;
wire u_usb_device_controller_usb_transact_inst_s_sendpid_3_17;
wire u_usb_device_controller_u_usb_packet_n640_22;
wire u_usb_device_controller_u_usb_packet_n640_23;
wire u_usb_device_controller_u_usb_packet_n642_22;
wire u_usb_device_controller_u_usb_packet_n642_23;
wire u_usb_device_controller_u_usb_packet_n644_22;
wire u_usb_device_controller_u_usb_packet_n644_23;
wire u_usb_device_controller_u_usb_packet_n646_21;
wire u_usb_device_controller_u_usb_packet_n646_22;
wire u_usb_device_controller_u_usb_packet_n646_23;
wire u_usb_device_controller_u_usb_packet_n650_22;
wire u_usb_device_controller_u_usb_packet_n650_23;
wire u_usb_device_controller_u_usb_packet_n650_24;
wire u_usb_device_controller_usb_control_inst_n1672_47;
wire u_usb_device_controller_usb_control_inst_n1672_48;
wire u_usb_device_controller_usb_control_inst_n1672_49;
wire u_usb_device_controller_usb_control_inst_n1680_48;
wire u_usb_device_controller_usb_control_inst_n1686_43;
wire u_usb_device_controller_usb_control_inst_n1686_44;
wire u_usb_device_controller_usb_control_inst_n1690_39;
wire u_usb_device_controller_u_usb_packet_n628_49;
wire u_usb_device_controller_u_usb_packet_n628_50;
wire u_usb_device_controller_u_usb_packet_n633_43;
wire u_usb_device_controller_u_usb_packet_n633_44;
wire u_usb_device_controller_usb_control_inst_n1860_33;
wire u_usb_device_controller_u_usb_init_n219_30;
wire u_usb_device_controller_n1534_35;
wire u_usb_device_controller_usbc_dsclen_0_20;
wire u_usb_device_controller_usbc_dsclen_0_21;
wire u_usb_device_controller_usbc_dsclen_0_22;
wire u_usb_device_controller_usbc_dsclen_0_23;
wire u_usb_device_controller_usbc_dsclen_1_21;
wire u_usb_device_controller_usbc_dsclen_1_22;
wire u_usb_device_controller_usbc_dsclen_2_18;
wire u_usb_device_controller_usbc_dsclen_2_19;
wire u_usb_device_controller_usbc_dsclen_2_20;
wire u_usb_device_controller_usbc_dsclen_3_18;
wire u_usb_device_controller_usbc_dsclen_3_19;
wire u_usb_device_controller_usbc_dsclen_3_20;
wire u_usb_device_controller_usbc_dsclen_4_19;
wire u_usb_device_controller_usbc_dsclen_5_18;
wire u_usb_device_controller_usbc_dsclen_5_19;
wire u_usb_device_controller_usbc_dsclen_5_20;
wire u_usb_device_controller_usbc_dsclen_6_18;
wire u_usb_device_controller_usbc_dsclen_6_19;
wire u_usb_device_controller_usbc_dsclen_6_20;
wire u_usb_device_controller_usbc_dsclen_7_18;
wire u_usb_device_controller_usbc_dsclen_7_19;
wire u_usb_device_controller_usbc_dsclen_7_20;
wire u_usb_device_controller_descrom_start_0_19;
wire u_usb_device_controller_descrom_start_1_19;
wire u_usb_device_controller_descrom_start_2_19;
wire u_usb_device_controller_descrom_start_3_19;
wire u_usb_device_controller_descrom_start_4_19;
wire u_usb_device_controller_descrom_start_5_19;
wire u_usb_device_controller_descrom_start_6_19;
wire u_usb_device_controller_descrom_start_7_19;
wire u_usb_device_controller_descrom_start_8_19;
wire u_usb_device_controller_descrom_start_9_19;
wire u_usb_device_controller_u_usb_packet_n771_13;
wire u_usb_device_controller_u_usb_packet_n771_14;
wire u_usb_device_controller_u_usb_packet_n767_9;
wire u_usb_device_controller_u_usb_packet_n767_10;
wire u_usb_device_controller_u_usb_packet_n912_22;
wire u_usb_device_controller_u_usb_packet_n912_23;
wire u_usb_device_controller_u_usb_init_n212_46;
wire u_usb_device_controller_u_usb_init_n212_47;
wire u_usb_device_controller_u_usb_init_n212_48;
wire u_usb_device_controller_u_usb_init_n212_49;
wire u_usb_device_controller_u_usb_init_n212_50;
wire u_usb_device_controller_u_usb_init_n212_51;
wire u_usb_device_controller_u_usb_init_n212_52;
wire u_usb_device_controller_u_usb_init_n212_53;
wire u_usb_device_controller_u_usb_init_n212_54;
wire u_usb_device_controller_u_usb_init_n215_61;
wire u_usb_device_controller_u_usb_init_n215_62;
wire u_usb_device_controller_u_usb_init_n215_63;
wire u_usb_device_controller_u_usb_packet_n328_25;
wire u_usb_device_controller_u_usb_init_s_state_3_16;
wire u_usb_device_controller_u_usb_init_s_chirpcnt_2_15;
wire u_usb_device_controller_u_usb_packet_n640_24;
wire u_usb_device_controller_u_usb_packet_n640_25;
wire u_usb_device_controller_u_usb_packet_n642_24;
wire u_usb_device_controller_u_usb_packet_n644_24;
wire u_usb_device_controller_u_usb_packet_n644_25;
wire u_usb_device_controller_u_usb_packet_n646_24;
wire u_usb_device_controller_u_usb_packet_n650_25;
wire u_usb_device_controller_usb_control_inst_n1860_34;
wire u_usb_device_controller_usbc_dsclen_0_24;
wire u_usb_device_controller_usbc_dsclen_6_21;
wire u_usb_device_controller_descrom_start_0_20;
wire u_usb_device_controller_descrom_start_1_20;
wire u_usb_device_controller_descrom_start_2_20;
wire u_usb_device_controller_descrom_start_3_20;
wire u_usb_device_controller_descrom_start_4_20;
wire u_usb_device_controller_descrom_start_5_20;
wire u_usb_device_controller_descrom_start_6_20;
wire u_usb_device_controller_descrom_start_7_20;
wire u_usb_device_controller_descrom_start_8_20;
wire u_usb_device_controller_descrom_start_9_20;
wire u_usb_device_controller_u_usb_packet_n771_15;
wire u_usb_device_controller_u_usb_packet_n771_16;
wire u_usb_device_controller_u_usb_init_n212_55;
wire u_usb_device_controller_usb_transact_inst_n1080_53;
wire u_usb_device_controller_n1266;
wire u_usb_device_controller_n1595_23;
wire u_usb_device_controller_n1601_23;
wire u_usb_device_controller_usb_control_inst_n1680_50;
wire u_usb_device_controller_utmi_dataout_o_d_7_10;
wire u_usb_device_controller_test_packet_inst_n315_10;
wire u_usb_device_controller_u_usb_init_n215_65;
wire u_usb_device_controller_u_usb_init_n212_57;
wire u_usb_device_controller_u_usb_init_n212_59;
wire u_usb_device_controller_u_usb_init_n215_67;
wire u_usb_device_controller_u_usb_init_n215_69;
wire u_usb_device_controller_u_usb_init_s_state_3_18;
wire u_usb_device_controller_u_usb_packet_crc5_buf_4_13;
wire u_usb_device_controller_u_usb_packet_n328_27;
wire u_usb_device_controller_u_usb_packet_n624;
wire u_usb_device_controller_u_usb_packet_n615_49;
wire u_usb_device_controller_u_usb_packet_n767_12;
wire u_usb_device_controller_u_usb_packet_n768;
wire u_usb_device_controller_u_usb_packet_n648;
wire u_usb_device_controller_u_usb_packet_n654;
wire u_usb_device_controller_usb_control_inst_n1655_18;
wire u_usb_device_controller_usb_control_inst_s_setupptr_2_12;
wire u_usb_device_controller_usb_control_inst_n1678_46;
wire u_usb_device_controller_usb_control_inst_n1761_16;
wire u_usb_device_controller_usb_control_inst_n1709_19;
wire u_usb_device_controller_usb_control_inst_n1909;
wire u_usb_device_controller_usb_transact_inst_n1099_49;
wire u_usb_device_controller_usb_transact_inst_s_sendpid_3;
wire u_usb_device_controller_usb_transact_inst_n1124_28;
wire u_usb_device_controller_usb_transact_inst_n1138_35;
wire u_usb_device_controller_usb_transact_inst_n1138_37;
wire u_usb_device_controller_usb_transact_inst_n1136_29;
wire u_usb_device_controller_usb_transact_inst_n1138_39;
wire u_usb_device_controller_usb_transact_inst_n1565;
wire u_usb_device_controller_usbc_dsclen_0;
wire u_usb_device_controller_usbc_dsclen_6;
wire u_usb_device_controller_n1607_23;
wire u_usb_device_controller_n1611;
wire u_usb_device_controller_n1810;
wire u_usb_device_controller_utmi_txvalid_o_d_6;
wire u_usb_device_controller_u_usb_init_n212_61;
wire u_usb_device_controller_u_usb_init_n212_63;
wire u_usb_device_controller_u_usb_init_n216_56;
wire u_usb_device_controller_u_usb_packet_n920_9;
wire u_usb_device_controller_u_usb_packet_PHY_TXVALID;
wire u_usb_device_controller_u_usb_packet_n1454;
wire u_usb_device_controller_u_usb_packet_n620;
wire u_usb_device_controller_usb_transact_inst_n1091_54;
wire u_usb_device_controller_u_usb_packet_n624_37;
wire u_usb_device_controller_u_usb_packet_n622_46;
wire u_usb_device_controller_u_usb_packet_n784_16;
wire u_usb_device_controller_u_usb_packet_n626_48;
wire u_usb_device_controller_usb_control_inst_n1686_48;
wire u_usb_device_controller_usb_control_inst_s_answerlen_7_11;
wire u_usb_device_controller_usb_control_inst_n2896_9;
wire u_usb_device_controller_usb_control_inst_n1661_22;
wire u_usb_device_controller_usb_control_inst_s_answerptr_5_14;
wire u_usb_device_controller_usb_control_inst_C_CLRIN_1_9;
wire u_usb_device_controller_usb_control_inst_s_interface_set;
wire u_usb_device_controller_usb_control_inst_s_answerlen_7_13;
wire u_usb_device_controller_usb_transact_inst_n1086_48;
wire u_usb_device_controller_usb_transact_inst_s_sendpid_3_21;
wire u_usb_device_controller_usb_transact_inst_n1142_25;
wire u_usb_device_controller_usb_transact_inst_n1148_25;
wire u_usb_device_controller_usb_transact_inst_n1086_50;
wire u_usb_device_controller_usb_transact_inst_n1138_41;
wire u_usb_device_controller_n1585;
wire u_usb_device_controller_n1529_31;
wire u_usb_device_controller_rxact_o_d;
wire u_usb_device_controller_test_packet_inst_n131_8;
wire u_usb_device_controller_test_packet_inst_n318_17;
wire u_usb_device_controller_u_usb_init_n210;
wire u_usb_device_controller_u_usb_init_n209;
wire u_usb_device_controller_u_usb_init_s_opmode_0;
wire u_usb_device_controller_u_usb_packet_n800_9;
wire u_usb_device_controller_u_usb_packet_n784_18;
wire u_usb_device_controller_usb_control_inst_n1649_23;
wire u_usb_device_controller_usb_control_inst_n1674;
wire u_usb_device_controller_descrom_start_0_23;
wire u_usb_device_controller_usb_control_inst_n1876_9;
wire u_usb_device_controller_usb_control_inst_n1836_13;
wire u_usb_device_controller_usb_control_inst_n1686_50;
wire u_usb_device_controller_usb_control_inst_n1693;
wire u_usb_device_controller_usb_control_inst_n2067;
wire u_usb_device_controller_usb_transact_inst_n1088_48;
wire u_usb_device_controller_usb_transact_inst_n1070_18;
wire u_usb_device_controller_usb_transact_inst_n1111;
wire u_usb_device_controller_usb_transact_inst_T_PING_7;
wire u_usb_device_controller_usb_transact_inst_n1041_8;
wire u_usb_device_controller_u_usb_packet_n770_10;
wire u_usb_device_controller_u_usb_packet_n770_12;
wire u_usb_device_controller_u_usb_packet_n640_27;
wire u_usb_device_controller_usb_transact_inst_txpop_o_d_9;
wire u_usb_device_controller_u_usb_init_s_state_2_18;
wire u_usb_device_controller_u_usb_init_n223;
wire u_usb_device_controller_u_usb_init_n214;
wire u_usb_device_controller_u_usb_init_s_chirpcnt_2;
wire u_usb_device_controller_u_usb_init_s_state_2_20;
wire u_usb_device_controller_u_usb_init_n212_65;
wire u_usb_device_controller_u_usb_init_n215_71;
wire u_usb_device_controller_u_usb_init_s_highspeed;
wire u_usb_device_controller_u_usb_init_n414;
wire u_usb_device_controller_u_usb_packet_crc16_buf_15_12;
wire u_usb_device_controller_usb_control_inst_n1701_21;
wire u_usb_device_controller_usb_control_inst_n1876_11;
wire u_usb_device_controller_usb_control_inst_n1864_8;
wire u_usb_device_controller_usb_control_inst_n1670_45;
wire u_usb_device_controller_usb_control_inst_n1836_15;
wire u_usb_device_controller_usb_transact_inst_n1080_55;
wire u_usb_device_controller_u_usb_packet_s_state_11_27;
wire u_usb_device_controller_n1240;
wire u_usb_device_controller_n503_10;
wire u_usb_device_controller_n443_10;
wire u_usb_device_controller_n385_10;
wire u_usb_device_controller_isync_3;
wire u_usb_device_controller_isync_2;
wire u_usb_device_controller_isync_1;
wire u_usb_device_controller_n1524_27;
wire u_usb_device_controller_n1534_37;
wire u_usb_device_controller_n384_10;
wire u_usb_device_controller_n1519_32;
wire u_usb_device_controller_n1520;
wire u_usb_device_controller_n1593_24;
wire u_usb_device_controller_setup_o_d;
wire u_usb_device_controller_test_packet_inst_n378_8;
wire u_usb_device_controller_usb_control_inst_n1876_13;
wire u_usb_device_controller_usb_control_inst_n1805;
wire u_usb_device_controller_usb_control_inst_n1775;
wire u_usb_device_controller_test_packet_inst_n312_13;
wire u_usb_device_controller_test_packet_inst_test_data_val_9;
wire u_usb_device_controller_usb_control_inst_n1773;
wire u_usb_device_controller_usb_control_inst_n1771;
wire u_usb_device_controller_usb_control_inst_n1769;
wire u_usb_device_controller_usb_control_inst_n1767;
wire u_usb_device_controller_usb_control_inst_n1765;
wire u_usb_device_controller_usb_control_inst_n1763;
wire u_usb_device_controller_usb_control_inst_n1761;
wire u_usb_device_controller_usb_control_inst_n1803;
wire u_usb_device_controller_usb_control_inst_n1801;
wire u_usb_device_controller_usb_control_inst_n1799;
wire u_usb_device_controller_usb_control_inst_n1797;
wire u_usb_device_controller_usb_control_inst_n1795;
wire u_usb_device_controller_usb_control_inst_n1793;
wire u_usb_device_controller_usb_control_inst_n1791;
wire u_usb_device_controller_usb_control_inst_n2902;
wire u_usb_device_controller_usb_control_inst_n1388_12;
wire u_usb_device_controller_usb_control_inst_n1676;
wire u_usb_device_controller_n1231_9;
wire u_usb_device_controller_n1167_9;
wire u_usb_device_controller_n1105_9;
wire u_usb_device_controller_n1043_9;
wire u_usb_device_controller_isync_15;
wire u_usb_device_controller_isync_14;
wire u_usb_device_controller_isync_13;
wire u_usb_device_controller_isync_12;
wire u_usb_device_controller_n743_9;
wire u_usb_device_controller_n681_9;
wire u_usb_device_controller_n621_9;
wire u_usb_device_controller_n561_10;
wire u_usb_device_controller_isync_7;
wire u_usb_device_controller_isync_6;
wire u_usb_device_controller_isync_5;
wire u_usb_device_controller_isync_4;
wire u_usb_device_controller_n983_9;
wire u_usb_device_controller_n921_9;
wire u_usb_device_controller_n861_9;
wire u_usb_device_controller_n801_9;
wire u_usb_device_controller_isync_11;
wire u_usb_device_controller_isync_10;
wire u_usb_device_controller_isync_9;
wire u_usb_device_controller_isync_8;
wire u_usb_device_controller_usb_control_inst_n1813;
wire u_usb_device_controller_usb_control_inst_n1783;
wire u_usb_device_controller_usb_control_inst_n1817;
wire u_usb_device_controller_usb_control_inst_n1787;
wire u_usb_device_controller_usb_control_inst_n1819;
wire u_usb_device_controller_usb_control_inst_n1789;
wire u_usb_device_controller_usb_control_inst_n1785;
wire u_usb_device_controller_usb_control_inst_n1781;
wire u_usb_device_controller_usb_control_inst_n1779;
wire u_usb_device_controller_usb_control_inst_n1777;
wire u_usb_device_controller_usb_control_inst_n1815;
wire u_usb_device_controller_usb_control_inst_n1811;
wire u_usb_device_controller_usb_control_inst_n1809;
wire u_usb_device_controller_usb_control_inst_n1807;
wire u_usb_device_controller_utmi_txvalid_o_d_8;
wire u_usb_device_controller_usb_control_inst_n1652_22;
wire u_usb_device_controller_usb_control_inst_s_sendbyte_7_19;
wire u_usb_device_controller_usb_transact_inst_n1101_48;
wire u_usb_device_controller_usb_transact_inst_n1070_20;
wire u_usb_device_controller_usb_transact_inst_n1076_24;
wire u_usb_device_controller_usb_transact_inst_n1163_24;
wire u_usb_device_controller_usb_transact_inst_n1068_16;
wire u_usb_device_controller_usb_transact_inst_n1076_26;
wire u_usb_device_controller_usb_transact_inst_n1064_23;
wire u_usb_device_controller_rxval_o_d;
wire u_usb_device_controller_n2393;
wire u_usb_device_controller_n1595;
wire u_usb_device_controller_n1601;
wire u_usb_device_controller_n1607;
wire u_usb_device_controller_n1613;
wire u_usb_device_controller_u_usb_packet_n328_29;
wire u_usb_device_controller_u_usb_packet_n328_31;
wire u_usb_device_controller_usbc_dsclen_1_24;
wire u_usb_device_controller_usbc_dsclen_1_26;
wire u_usb_device_controller_usbc_dsclen_0_28;
wire u_usb_device_controller_usb_transact_inst_n1068_18;
wire u_usb_device_controller_u_usb_packet_crc16_buf_15_14;
wire u_usb_device_controller_usb_transact_inst_n1086_52;
wire u_usb_device_controller_usb_transact_inst_n1111_22;
wire u_usb_device_controller_usb_transact_inst_s_endpt_0_9;
wire u_usb_device_controller_n2393_9;
wire u_usb_device_controller_usb_transact_inst_s_endpt_3;
wire u_usb_device_controller_u_usb_packet_n773;
wire u_usb_device_controller_u_usb_packet_n769;
wire u_usb_device_controller_u_usb_packet_n772;
wire u_usb_device_controller_u_usb_packet_n762;
wire u_usb_device_controller_u_usb_packet_n763;
wire u_usb_device_controller_u_usb_packet_n765;
wire u_usb_device_controller_u_usb_packet_n766;
wire u_usb_device_controller_u_usb_packet_n767;
wire u_usb_device_controller_u_usb_packet_n770;
wire u_usb_device_controller_u_usb_packet_n771;
wire u_usb_device_controller_u_usb_packet_n774;
wire u_usb_device_controller_u_usb_packet_n784_20;
wire u_usb_device_controller_u_usb_init_s_state_2;
wire u_usb_device_controller_usb_control_inst_n1652_24;
wire u_usb_device_controller_usb_control_inst_s_sendbyte_7;
wire u_usb_device_controller_usb_transact_inst_n1091_56;
wire u_usb_device_controller_usb_transact_inst_n1140;
wire u_usb_device_controller_usb_transact_inst_s_sendpid_3_23;
wire u_usb_device_controller_u_usb_packet_n622;
wire u_usb_device_controller_usb_transact_inst_n1107_48;
wire u_usb_device_controller_usb_transact_inst_n1064_25;
wire u_usb_device_controller_usb_transact_inst_s_endpt_0;
wire u_usb_device_controller_usb_control_inst_n1674_44;
wire u_usb_device_controller_usb_control_inst_s_ctlparam_7;
wire u_usb_device_controller_usb_transact_inst_n1099;
wire u_usb_device_controller_usb_transact_inst_wait_count_9;
wire u_usb_device_controller_s_bufptr_1;
wire u_usb_device_controller_usb_control_inst_usbc_dscrd;
wire u_usb_device_controller_usb_transact_inst_n1064_27;
wire u_usb_device_controller_usb_transact_inst_n1138_43;
wire u_usb_device_controller_n1716;
wire u_usb_device_controller_n1714;
wire u_usb_device_controller_n1713;
wire u_usb_device_controller_n1712;
wire u_usb_device_controller_n1711;
wire u_usb_device_controller_n1710;
wire u_usb_device_controller_n1709;
wire u_usb_device_controller_n1708;
wire u_usb_device_controller_n1707;
wire u_usb_device_controller_n1706;
wire u_usb_device_controller_n1705;
wire u_usb_device_controller_n1704;
wire u_usb_device_controller_n1703;
wire u_usb_device_controller_n1702;
wire u_usb_device_controller_n1701;
wire u_usb_device_controller_n1700;
wire u_usb_device_controller_n1699;
wire u_usb_device_controller_n1760;
wire u_usb_device_controller_n1761;
wire u_usb_device_controller_n1762;
wire u_usb_device_controller_n1763;
wire u_usb_device_controller_n1764;
wire u_usb_device_controller_n1765;
wire u_usb_device_controller_n1766;
wire u_usb_device_controller_n1767;
wire u_usb_device_controller_n1770;
wire u_usb_device_controller_u_usb_init_n241;
wire u_usb_device_controller_u_usb_init_n279;
wire u_usb_device_controller_usb_control_inst_n1699_15;
wire u_usb_device_controller_usb_control_inst_n1699;
wire u_usb_device_controller_usb_control_inst_s_setupptr_2;
wire u_usb_device_controller_n340;
wire u_usb_device_controller_n395;
wire u_usb_device_controller_n398;
wire u_usb_device_controller_n453;
wire u_usb_device_controller_n456;
wire u_usb_device_controller_n513;
wire u_usb_device_controller_n516;
wire u_usb_device_controller_n571;
wire u_usb_device_controller_n574;
wire u_usb_device_controller_n631;
wire u_usb_device_controller_n634;
wire u_usb_device_controller_n691;
wire u_usb_device_controller_n694;
wire u_usb_device_controller_n753;
wire u_usb_device_controller_n756;
wire u_usb_device_controller_n811;
wire u_usb_device_controller_n814;
wire u_usb_device_controller_n871;
wire u_usb_device_controller_n874;
wire u_usb_device_controller_n931;
wire u_usb_device_controller_n934;
wire u_usb_device_controller_n993;
wire u_usb_device_controller_n996;
wire u_usb_device_controller_n1053;
wire u_usb_device_controller_n1056;
wire u_usb_device_controller_n1115;
wire u_usb_device_controller_n1118;
wire u_usb_device_controller_n1177;
wire u_usb_device_controller_n1180;
wire u_usb_device_controller_n337;
wire u_usb_device_controller_n2024;
wire u_usb_device_controller_n2024_11;
wire u_usb_device_controller_u_usb_init_n316;
wire GND;
wire VCC;
wire [9:0] desc_dev_addr_i_d;
wire [7:0] desc_dev_len_i_d;
wire [9:0] desc_fscfg_addr_i_d;
wire [7:0] desc_fscfg_len_i_d;
wire [9:0] desc_hscfg_addr_i_d;
wire [7:0] desc_hscfg_len_i_d;
wire [9:0] desc_oscfg_addr_i_d;
wire [9:0] desc_qual_addr_i_d;
wire [7:0] desc_qual_len_i_d;
wire [9:0] desc_strlang_addr_i_d;
wire [9:0] desc_strproduct_addr_i_d;
wire [7:0] desc_strproduct_len_i_d;
wire [9:0] desc_strserial_addr_i_d;
wire [7:0] desc_strserial_len_i_d;
wire [9:0] desc_strvendor_addr_i_d;
wire [7:0] desc_strvendor_len_i_d;
wire [7:0] descrom_rdata_i_d;
wire [7:0] inf_alter_i_d;
wire [7:0] txdat_i_d;
wire [11:0] txdat_len_i_d;
wire [3:0] u_usb_device_controller_cur_state;
wire [9:0] u_usb_device_controller_descrom_raddr_o_d;
wire [15:1] u_usb_device_controller_halt_in;
wire [15:1] u_usb_device_controller_halt_out;
wire [15:1] u_usb_device_controller_isync;
wire [3:0] u_usb_device_controller_next_state;
wire [15:1] u_usb_device_controller_osync;
wire [7:0] u_usb_device_controller_rxdat_d0;
wire [7:0] u_usb_device_controller_rxdat_d1;
wire [7:0] u_usb_device_controller_rxdat_d2;
wire [7:0] u_usb_device_controller_rxdat_o_d;
wire [11:0] u_usb_device_controller_s_bufptr;
wire [11:0] u_usb_device_controller_s_txbuf_stop;
wire [11:0] u_usb_device_controller_test_packet_inst_cnt;
wire [7:0] u_usb_device_controller_test_packet_inst_test_data_Z;
wire [2:0] u_usb_device_controller_u_usb_init_s_chirpcnt;
wire [1:0] u_usb_device_controller_u_usb_init_s_linestate;
wire [3:1] u_usb_device_controller_u_usb_init_s_state;
wire [15:0] u_usb_device_controller_u_usb_init_s_timer1;
wire [19:0] u_usb_device_controller_u_usb_init_s_timer2;
wire [0:0] u_usb_device_controller_u_usb_init_s_usb_test_en;
wire [1:0] u_usb_device_controller_u_usb_init_usbi_opmode;
wire [0:0] u_usb_device_controller_u_usb_init_utmi_xcvrselect_o_d;
wire [15:0] u_usb_device_controller_u_usb_packet_crc16_buf;
wire [4:0] u_usb_device_controller_u_usb_packet_crc5_buf;
wire [7:0] u_usb_device_controller_u_usb_packet_s_dataout;
wire [8:0] u_usb_device_controller_u_usb_packet_s_state;
wire [7:0] u_usb_device_controller_u_usb_packet_usbp_dataout_o;
wire [7:0] u_usb_device_controller_u_usb_packet_usbt_rxdat;
wire [7:0] u_usb_device_controller_usb_control_inst_inf_alter_o_d;
wire [7:0] u_usb_device_controller_usb_control_inst_inf_sel_o_d;
wire [7:0] u_usb_device_controller_usb_control_inst_s_answerlen;
wire [3:0] u_usb_device_controller_usb_control_inst_s_ctlrequest;
wire [2:0] u_usb_device_controller_usb_control_inst_s_setupptr;
wire [9:0] u_usb_device_controller_usb_control_inst_s_state;
wire [6:0] u_usb_device_controller_usb_control_inst_usbc_addr;
wire [15:1] u_usb_device_controller_usb_control_inst_usbc_clr_in;
wire [15:1] u_usb_device_controller_usb_control_inst_usbc_clr_out;
wire [7:0] u_usb_device_controller_usb_control_inst_usbc_dscinx;
wire [7:0] u_usb_device_controller_usb_control_inst_usbc_dscoff;
wire [2:0] u_usb_device_controller_usb_control_inst_usbc_dsctyp;
wire [15:1] u_usb_device_controller_usb_control_inst_usbc_sethlt_in;
wire [15:1] u_usb_device_controller_usb_control_inst_usbc_sethlt_out;
wire [7:0] u_usb_device_controller_usb_control_inst_usbc_testmode;
wire [7:0] u_usb_device_controller_usb_control_inst_usbc_txdat;
wire [3:0] u_usb_device_controller_usb_transact_inst_endpt_o_d;
wire [3:0] u_usb_device_controller_usb_transact_inst_s_sendpid;
wire [12:0] u_usb_device_controller_usb_transact_inst_s_state;
wire [15:0] u_usb_device_controller_usb_transact_inst_wait_count;
wire [7:0] u_usb_device_controller_utmi_dataout_o_d;
wire [1:0] u_usb_device_controller_utmi_opmode_o_d;
wire [7:0] utmi_datain_i_d;
wire [1:0] utmi_linestate_i_d;
  IBUF clk_i_ibuf (
    .O(clk_i_d),
    .I(clk_i) 
);
  IBUF reset_i_ibuf (
    .O(reset_i_d),
    .I(reset_i) 
);
  IBUF txdat_i_0_ibuf (
    .O(txdat_i_d[0]),
    .I(txdat_i[0]) 
);
  IBUF txdat_i_1_ibuf (
    .O(txdat_i_d[1]),
    .I(txdat_i[1]) 
);
  IBUF txdat_i_2_ibuf (
    .O(txdat_i_d[2]),
    .I(txdat_i[2]) 
);
  IBUF txdat_i_3_ibuf (
    .O(txdat_i_d[3]),
    .I(txdat_i[3]) 
);
  IBUF txdat_i_4_ibuf (
    .O(txdat_i_d[4]),
    .I(txdat_i[4]) 
);
  IBUF txdat_i_5_ibuf (
    .O(txdat_i_d[5]),
    .I(txdat_i[5]) 
);
  IBUF txdat_i_6_ibuf (
    .O(txdat_i_d[6]),
    .I(txdat_i[6]) 
);
  IBUF txdat_i_7_ibuf (
    .O(txdat_i_d[7]),
    .I(txdat_i[7]) 
);
  IBUF txval_i_ibuf (
    .O(txval_i_d),
    .I(txval_i) 
);
  IBUF txdat_len_i_0_ibuf (
    .O(txdat_len_i_d[0]),
    .I(txdat_len_i[0]) 
);
  IBUF txdat_len_i_1_ibuf (
    .O(txdat_len_i_d[1]),
    .I(txdat_len_i[1]) 
);
  IBUF txdat_len_i_2_ibuf (
    .O(txdat_len_i_d[2]),
    .I(txdat_len_i[2]) 
);
  IBUF txdat_len_i_3_ibuf (
    .O(txdat_len_i_d[3]),
    .I(txdat_len_i[3]) 
);
  IBUF txdat_len_i_4_ibuf (
    .O(txdat_len_i_d[4]),
    .I(txdat_len_i[4]) 
);
  IBUF txdat_len_i_5_ibuf (
    .O(txdat_len_i_d[5]),
    .I(txdat_len_i[5]) 
);
  IBUF txdat_len_i_6_ibuf (
    .O(txdat_len_i_d[6]),
    .I(txdat_len_i[6]) 
);
  IBUF txdat_len_i_7_ibuf (
    .O(txdat_len_i_d[7]),
    .I(txdat_len_i[7]) 
);
  IBUF txdat_len_i_8_ibuf (
    .O(txdat_len_i_d[8]),
    .I(txdat_len_i[8]) 
);
  IBUF txdat_len_i_9_ibuf (
    .O(txdat_len_i_d[9]),
    .I(txdat_len_i[9]) 
);
  IBUF txdat_len_i_10_ibuf (
    .O(txdat_len_i_d[10]),
    .I(txdat_len_i[10]) 
);
  IBUF txdat_len_i_11_ibuf (
    .O(txdat_len_i_d[11]),
    .I(txdat_len_i[11]) 
);
  IBUF txcork_i_ibuf (
    .O(txcork_i_d),
    .I(txcork_i) 
);
  IBUF rxrdy_i_ibuf (
    .O(rxrdy_i_d),
    .I(rxrdy_i) 
);
  IBUF inf_alter_i_0_ibuf (
    .O(inf_alter_i_d[0]),
    .I(inf_alter_i[0]) 
);
  IBUF inf_alter_i_1_ibuf (
    .O(inf_alter_i_d[1]),
    .I(inf_alter_i[1]) 
);
  IBUF inf_alter_i_2_ibuf (
    .O(inf_alter_i_d[2]),
    .I(inf_alter_i[2]) 
);
  IBUF inf_alter_i_3_ibuf (
    .O(inf_alter_i_d[3]),
    .I(inf_alter_i[3]) 
);
  IBUF inf_alter_i_4_ibuf (
    .O(inf_alter_i_d[4]),
    .I(inf_alter_i[4]) 
);
  IBUF inf_alter_i_5_ibuf (
    .O(inf_alter_i_d[5]),
    .I(inf_alter_i[5]) 
);
  IBUF inf_alter_i_6_ibuf (
    .O(inf_alter_i_d[6]),
    .I(inf_alter_i[6]) 
);
  IBUF inf_alter_i_7_ibuf (
    .O(inf_alter_i_d[7]),
    .I(inf_alter_i[7]) 
);
  IBUF descrom_rdata_i_0_ibuf (
    .O(descrom_rdata_i_d[0]),
    .I(descrom_rdata_i[0]) 
);
  IBUF descrom_rdata_i_1_ibuf (
    .O(descrom_rdata_i_d[1]),
    .I(descrom_rdata_i[1]) 
);
  IBUF descrom_rdata_i_2_ibuf (
    .O(descrom_rdata_i_d[2]),
    .I(descrom_rdata_i[2]) 
);
  IBUF descrom_rdata_i_3_ibuf (
    .O(descrom_rdata_i_d[3]),
    .I(descrom_rdata_i[3]) 
);
  IBUF descrom_rdata_i_4_ibuf (
    .O(descrom_rdata_i_d[4]),
    .I(descrom_rdata_i[4]) 
);
  IBUF descrom_rdata_i_5_ibuf (
    .O(descrom_rdata_i_d[5]),
    .I(descrom_rdata_i[5]) 
);
  IBUF descrom_rdata_i_6_ibuf (
    .O(descrom_rdata_i_d[6]),
    .I(descrom_rdata_i[6]) 
);
  IBUF descrom_rdata_i_7_ibuf (
    .O(descrom_rdata_i_d[7]),
    .I(descrom_rdata_i[7]) 
);
  IBUF desc_dev_addr_i_0_ibuf (
    .O(desc_dev_addr_i_d[0]),
    .I(desc_dev_addr_i[0]) 
);
  IBUF desc_dev_addr_i_1_ibuf (
    .O(desc_dev_addr_i_d[1]),
    .I(desc_dev_addr_i[1]) 
);
  IBUF desc_dev_addr_i_2_ibuf (
    .O(desc_dev_addr_i_d[2]),
    .I(desc_dev_addr_i[2]) 
);
  IBUF desc_dev_addr_i_3_ibuf (
    .O(desc_dev_addr_i_d[3]),
    .I(desc_dev_addr_i[3]) 
);
  IBUF desc_dev_addr_i_4_ibuf (
    .O(desc_dev_addr_i_d[4]),
    .I(desc_dev_addr_i[4]) 
);
  IBUF desc_dev_addr_i_5_ibuf (
    .O(desc_dev_addr_i_d[5]),
    .I(desc_dev_addr_i[5]) 
);
  IBUF desc_dev_addr_i_6_ibuf (
    .O(desc_dev_addr_i_d[6]),
    .I(desc_dev_addr_i[6]) 
);
  IBUF desc_dev_addr_i_7_ibuf (
    .O(desc_dev_addr_i_d[7]),
    .I(desc_dev_addr_i[7]) 
);
  IBUF desc_dev_addr_i_8_ibuf (
    .O(desc_dev_addr_i_d[8]),
    .I(desc_dev_addr_i[8]) 
);
  IBUF desc_dev_addr_i_9_ibuf (
    .O(desc_dev_addr_i_d[9]),
    .I(desc_dev_addr_i[9]) 
);
  IBUF desc_dev_len_i_0_ibuf (
    .O(desc_dev_len_i_d[0]),
    .I(desc_dev_len_i[0]) 
);
  IBUF desc_dev_len_i_1_ibuf (
    .O(desc_dev_len_i_d[1]),
    .I(desc_dev_len_i[1]) 
);
  IBUF desc_dev_len_i_2_ibuf (
    .O(desc_dev_len_i_d[2]),
    .I(desc_dev_len_i[2]) 
);
  IBUF desc_dev_len_i_3_ibuf (
    .O(desc_dev_len_i_d[3]),
    .I(desc_dev_len_i[3]) 
);
  IBUF desc_dev_len_i_4_ibuf (
    .O(desc_dev_len_i_d[4]),
    .I(desc_dev_len_i[4]) 
);
  IBUF desc_dev_len_i_5_ibuf (
    .O(desc_dev_len_i_d[5]),
    .I(desc_dev_len_i[5]) 
);
  IBUF desc_dev_len_i_6_ibuf (
    .O(desc_dev_len_i_d[6]),
    .I(desc_dev_len_i[6]) 
);
  IBUF desc_dev_len_i_7_ibuf (
    .O(desc_dev_len_i_d[7]),
    .I(desc_dev_len_i[7]) 
);
  IBUF desc_qual_addr_i_0_ibuf (
    .O(desc_qual_addr_i_d[0]),
    .I(desc_qual_addr_i[0]) 
);
  IBUF desc_qual_addr_i_1_ibuf (
    .O(desc_qual_addr_i_d[1]),
    .I(desc_qual_addr_i[1]) 
);
  IBUF desc_qual_addr_i_2_ibuf (
    .O(desc_qual_addr_i_d[2]),
    .I(desc_qual_addr_i[2]) 
);
  IBUF desc_qual_addr_i_3_ibuf (
    .O(desc_qual_addr_i_d[3]),
    .I(desc_qual_addr_i[3]) 
);
  IBUF desc_qual_addr_i_4_ibuf (
    .O(desc_qual_addr_i_d[4]),
    .I(desc_qual_addr_i[4]) 
);
  IBUF desc_qual_addr_i_5_ibuf (
    .O(desc_qual_addr_i_d[5]),
    .I(desc_qual_addr_i[5]) 
);
  IBUF desc_qual_addr_i_6_ibuf (
    .O(desc_qual_addr_i_d[6]),
    .I(desc_qual_addr_i[6]) 
);
  IBUF desc_qual_addr_i_7_ibuf (
    .O(desc_qual_addr_i_d[7]),
    .I(desc_qual_addr_i[7]) 
);
  IBUF desc_qual_addr_i_8_ibuf (
    .O(desc_qual_addr_i_d[8]),
    .I(desc_qual_addr_i[8]) 
);
  IBUF desc_qual_addr_i_9_ibuf (
    .O(desc_qual_addr_i_d[9]),
    .I(desc_qual_addr_i[9]) 
);
  IBUF desc_qual_len_i_0_ibuf (
    .O(desc_qual_len_i_d[0]),
    .I(desc_qual_len_i[0]) 
);
  IBUF desc_qual_len_i_1_ibuf (
    .O(desc_qual_len_i_d[1]),
    .I(desc_qual_len_i[1]) 
);
  IBUF desc_qual_len_i_2_ibuf (
    .O(desc_qual_len_i_d[2]),
    .I(desc_qual_len_i[2]) 
);
  IBUF desc_qual_len_i_3_ibuf (
    .O(desc_qual_len_i_d[3]),
    .I(desc_qual_len_i[3]) 
);
  IBUF desc_qual_len_i_4_ibuf (
    .O(desc_qual_len_i_d[4]),
    .I(desc_qual_len_i[4]) 
);
  IBUF desc_qual_len_i_5_ibuf (
    .O(desc_qual_len_i_d[5]),
    .I(desc_qual_len_i[5]) 
);
  IBUF desc_qual_len_i_6_ibuf (
    .O(desc_qual_len_i_d[6]),
    .I(desc_qual_len_i[6]) 
);
  IBUF desc_qual_len_i_7_ibuf (
    .O(desc_qual_len_i_d[7]),
    .I(desc_qual_len_i[7]) 
);
  IBUF desc_fscfg_addr_i_0_ibuf (
    .O(desc_fscfg_addr_i_d[0]),
    .I(desc_fscfg_addr_i[0]) 
);
  IBUF desc_fscfg_addr_i_1_ibuf (
    .O(desc_fscfg_addr_i_d[1]),
    .I(desc_fscfg_addr_i[1]) 
);
  IBUF desc_fscfg_addr_i_2_ibuf (
    .O(desc_fscfg_addr_i_d[2]),
    .I(desc_fscfg_addr_i[2]) 
);
  IBUF desc_fscfg_addr_i_3_ibuf (
    .O(desc_fscfg_addr_i_d[3]),
    .I(desc_fscfg_addr_i[3]) 
);
  IBUF desc_fscfg_addr_i_4_ibuf (
    .O(desc_fscfg_addr_i_d[4]),
    .I(desc_fscfg_addr_i[4]) 
);
  IBUF desc_fscfg_addr_i_5_ibuf (
    .O(desc_fscfg_addr_i_d[5]),
    .I(desc_fscfg_addr_i[5]) 
);
  IBUF desc_fscfg_addr_i_6_ibuf (
    .O(desc_fscfg_addr_i_d[6]),
    .I(desc_fscfg_addr_i[6]) 
);
  IBUF desc_fscfg_addr_i_7_ibuf (
    .O(desc_fscfg_addr_i_d[7]),
    .I(desc_fscfg_addr_i[7]) 
);
  IBUF desc_fscfg_addr_i_8_ibuf (
    .O(desc_fscfg_addr_i_d[8]),
    .I(desc_fscfg_addr_i[8]) 
);
  IBUF desc_fscfg_addr_i_9_ibuf (
    .O(desc_fscfg_addr_i_d[9]),
    .I(desc_fscfg_addr_i[9]) 
);
  IBUF desc_fscfg_len_i_0_ibuf (
    .O(desc_fscfg_len_i_d[0]),
    .I(desc_fscfg_len_i[0]) 
);
  IBUF desc_fscfg_len_i_1_ibuf (
    .O(desc_fscfg_len_i_d[1]),
    .I(desc_fscfg_len_i[1]) 
);
  IBUF desc_fscfg_len_i_2_ibuf (
    .O(desc_fscfg_len_i_d[2]),
    .I(desc_fscfg_len_i[2]) 
);
  IBUF desc_fscfg_len_i_3_ibuf (
    .O(desc_fscfg_len_i_d[3]),
    .I(desc_fscfg_len_i[3]) 
);
  IBUF desc_fscfg_len_i_4_ibuf (
    .O(desc_fscfg_len_i_d[4]),
    .I(desc_fscfg_len_i[4]) 
);
  IBUF desc_fscfg_len_i_5_ibuf (
    .O(desc_fscfg_len_i_d[5]),
    .I(desc_fscfg_len_i[5]) 
);
  IBUF desc_fscfg_len_i_6_ibuf (
    .O(desc_fscfg_len_i_d[6]),
    .I(desc_fscfg_len_i[6]) 
);
  IBUF desc_fscfg_len_i_7_ibuf (
    .O(desc_fscfg_len_i_d[7]),
    .I(desc_fscfg_len_i[7]) 
);
  IBUF desc_hscfg_addr_i_0_ibuf (
    .O(desc_hscfg_addr_i_d[0]),
    .I(desc_hscfg_addr_i[0]) 
);
  IBUF desc_hscfg_addr_i_1_ibuf (
    .O(desc_hscfg_addr_i_d[1]),
    .I(desc_hscfg_addr_i[1]) 
);
  IBUF desc_hscfg_addr_i_2_ibuf (
    .O(desc_hscfg_addr_i_d[2]),
    .I(desc_hscfg_addr_i[2]) 
);
  IBUF desc_hscfg_addr_i_3_ibuf (
    .O(desc_hscfg_addr_i_d[3]),
    .I(desc_hscfg_addr_i[3]) 
);
  IBUF desc_hscfg_addr_i_4_ibuf (
    .O(desc_hscfg_addr_i_d[4]),
    .I(desc_hscfg_addr_i[4]) 
);
  IBUF desc_hscfg_addr_i_5_ibuf (
    .O(desc_hscfg_addr_i_d[5]),
    .I(desc_hscfg_addr_i[5]) 
);
  IBUF desc_hscfg_addr_i_6_ibuf (
    .O(desc_hscfg_addr_i_d[6]),
    .I(desc_hscfg_addr_i[6]) 
);
  IBUF desc_hscfg_addr_i_7_ibuf (
    .O(desc_hscfg_addr_i_d[7]),
    .I(desc_hscfg_addr_i[7]) 
);
  IBUF desc_hscfg_addr_i_8_ibuf (
    .O(desc_hscfg_addr_i_d[8]),
    .I(desc_hscfg_addr_i[8]) 
);
  IBUF desc_hscfg_addr_i_9_ibuf (
    .O(desc_hscfg_addr_i_d[9]),
    .I(desc_hscfg_addr_i[9]) 
);
  IBUF desc_hscfg_len_i_0_ibuf (
    .O(desc_hscfg_len_i_d[0]),
    .I(desc_hscfg_len_i[0]) 
);
  IBUF desc_hscfg_len_i_1_ibuf (
    .O(desc_hscfg_len_i_d[1]),
    .I(desc_hscfg_len_i[1]) 
);
  IBUF desc_hscfg_len_i_2_ibuf (
    .O(desc_hscfg_len_i_d[2]),
    .I(desc_hscfg_len_i[2]) 
);
  IBUF desc_hscfg_len_i_3_ibuf (
    .O(desc_hscfg_len_i_d[3]),
    .I(desc_hscfg_len_i[3]) 
);
  IBUF desc_hscfg_len_i_4_ibuf (
    .O(desc_hscfg_len_i_d[4]),
    .I(desc_hscfg_len_i[4]) 
);
  IBUF desc_hscfg_len_i_5_ibuf (
    .O(desc_hscfg_len_i_d[5]),
    .I(desc_hscfg_len_i[5]) 
);
  IBUF desc_hscfg_len_i_6_ibuf (
    .O(desc_hscfg_len_i_d[6]),
    .I(desc_hscfg_len_i[6]) 
);
  IBUF desc_hscfg_len_i_7_ibuf (
    .O(desc_hscfg_len_i_d[7]),
    .I(desc_hscfg_len_i[7]) 
);
  IBUF desc_oscfg_addr_i_0_ibuf (
    .O(desc_oscfg_addr_i_d[0]),
    .I(desc_oscfg_addr_i[0]) 
);
  IBUF desc_oscfg_addr_i_1_ibuf (
    .O(desc_oscfg_addr_i_d[1]),
    .I(desc_oscfg_addr_i[1]) 
);
  IBUF desc_oscfg_addr_i_2_ibuf (
    .O(desc_oscfg_addr_i_d[2]),
    .I(desc_oscfg_addr_i[2]) 
);
  IBUF desc_oscfg_addr_i_3_ibuf (
    .O(desc_oscfg_addr_i_d[3]),
    .I(desc_oscfg_addr_i[3]) 
);
  IBUF desc_oscfg_addr_i_4_ibuf (
    .O(desc_oscfg_addr_i_d[4]),
    .I(desc_oscfg_addr_i[4]) 
);
  IBUF desc_oscfg_addr_i_5_ibuf (
    .O(desc_oscfg_addr_i_d[5]),
    .I(desc_oscfg_addr_i[5]) 
);
  IBUF desc_oscfg_addr_i_6_ibuf (
    .O(desc_oscfg_addr_i_d[6]),
    .I(desc_oscfg_addr_i[6]) 
);
  IBUF desc_oscfg_addr_i_7_ibuf (
    .O(desc_oscfg_addr_i_d[7]),
    .I(desc_oscfg_addr_i[7]) 
);
  IBUF desc_oscfg_addr_i_8_ibuf (
    .O(desc_oscfg_addr_i_d[8]),
    .I(desc_oscfg_addr_i[8]) 
);
  IBUF desc_oscfg_addr_i_9_ibuf (
    .O(desc_oscfg_addr_i_d[9]),
    .I(desc_oscfg_addr_i[9]) 
);
  IBUF desc_strlang_addr_i_0_ibuf (
    .O(desc_strlang_addr_i_d[0]),
    .I(desc_strlang_addr_i[0]) 
);
  IBUF desc_strlang_addr_i_1_ibuf (
    .O(desc_strlang_addr_i_d[1]),
    .I(desc_strlang_addr_i[1]) 
);
  IBUF desc_strlang_addr_i_2_ibuf (
    .O(desc_strlang_addr_i_d[2]),
    .I(desc_strlang_addr_i[2]) 
);
  IBUF desc_strlang_addr_i_3_ibuf (
    .O(desc_strlang_addr_i_d[3]),
    .I(desc_strlang_addr_i[3]) 
);
  IBUF desc_strlang_addr_i_4_ibuf (
    .O(desc_strlang_addr_i_d[4]),
    .I(desc_strlang_addr_i[4]) 
);
  IBUF desc_strlang_addr_i_5_ibuf (
    .O(desc_strlang_addr_i_d[5]),
    .I(desc_strlang_addr_i[5]) 
);
  IBUF desc_strlang_addr_i_6_ibuf (
    .O(desc_strlang_addr_i_d[6]),
    .I(desc_strlang_addr_i[6]) 
);
  IBUF desc_strlang_addr_i_7_ibuf (
    .O(desc_strlang_addr_i_d[7]),
    .I(desc_strlang_addr_i[7]) 
);
  IBUF desc_strlang_addr_i_8_ibuf (
    .O(desc_strlang_addr_i_d[8]),
    .I(desc_strlang_addr_i[8]) 
);
  IBUF desc_strlang_addr_i_9_ibuf (
    .O(desc_strlang_addr_i_d[9]),
    .I(desc_strlang_addr_i[9]) 
);
  IBUF desc_strvendor_addr_i_0_ibuf (
    .O(desc_strvendor_addr_i_d[0]),
    .I(desc_strvendor_addr_i[0]) 
);
  IBUF desc_strvendor_addr_i_1_ibuf (
    .O(desc_strvendor_addr_i_d[1]),
    .I(desc_strvendor_addr_i[1]) 
);
  IBUF desc_strvendor_addr_i_2_ibuf (
    .O(desc_strvendor_addr_i_d[2]),
    .I(desc_strvendor_addr_i[2]) 
);
  IBUF desc_strvendor_addr_i_3_ibuf (
    .O(desc_strvendor_addr_i_d[3]),
    .I(desc_strvendor_addr_i[3]) 
);
  IBUF desc_strvendor_addr_i_4_ibuf (
    .O(desc_strvendor_addr_i_d[4]),
    .I(desc_strvendor_addr_i[4]) 
);
  IBUF desc_strvendor_addr_i_5_ibuf (
    .O(desc_strvendor_addr_i_d[5]),
    .I(desc_strvendor_addr_i[5]) 
);
  IBUF desc_strvendor_addr_i_6_ibuf (
    .O(desc_strvendor_addr_i_d[6]),
    .I(desc_strvendor_addr_i[6]) 
);
  IBUF desc_strvendor_addr_i_7_ibuf (
    .O(desc_strvendor_addr_i_d[7]),
    .I(desc_strvendor_addr_i[7]) 
);
  IBUF desc_strvendor_addr_i_8_ibuf (
    .O(desc_strvendor_addr_i_d[8]),
    .I(desc_strvendor_addr_i[8]) 
);
  IBUF desc_strvendor_addr_i_9_ibuf (
    .O(desc_strvendor_addr_i_d[9]),
    .I(desc_strvendor_addr_i[9]) 
);
  IBUF desc_strvendor_len_i_0_ibuf (
    .O(desc_strvendor_len_i_d[0]),
    .I(desc_strvendor_len_i[0]) 
);
  IBUF desc_strvendor_len_i_1_ibuf (
    .O(desc_strvendor_len_i_d[1]),
    .I(desc_strvendor_len_i[1]) 
);
  IBUF desc_strvendor_len_i_2_ibuf (
    .O(desc_strvendor_len_i_d[2]),
    .I(desc_strvendor_len_i[2]) 
);
  IBUF desc_strvendor_len_i_3_ibuf (
    .O(desc_strvendor_len_i_d[3]),
    .I(desc_strvendor_len_i[3]) 
);
  IBUF desc_strvendor_len_i_4_ibuf (
    .O(desc_strvendor_len_i_d[4]),
    .I(desc_strvendor_len_i[4]) 
);
  IBUF desc_strvendor_len_i_5_ibuf (
    .O(desc_strvendor_len_i_d[5]),
    .I(desc_strvendor_len_i[5]) 
);
  IBUF desc_strvendor_len_i_6_ibuf (
    .O(desc_strvendor_len_i_d[6]),
    .I(desc_strvendor_len_i[6]) 
);
  IBUF desc_strvendor_len_i_7_ibuf (
    .O(desc_strvendor_len_i_d[7]),
    .I(desc_strvendor_len_i[7]) 
);
  IBUF desc_strproduct_addr_i_0_ibuf (
    .O(desc_strproduct_addr_i_d[0]),
    .I(desc_strproduct_addr_i[0]) 
);
  IBUF desc_strproduct_addr_i_1_ibuf (
    .O(desc_strproduct_addr_i_d[1]),
    .I(desc_strproduct_addr_i[1]) 
);
  IBUF desc_strproduct_addr_i_2_ibuf (
    .O(desc_strproduct_addr_i_d[2]),
    .I(desc_strproduct_addr_i[2]) 
);
  IBUF desc_strproduct_addr_i_3_ibuf (
    .O(desc_strproduct_addr_i_d[3]),
    .I(desc_strproduct_addr_i[3]) 
);
  IBUF desc_strproduct_addr_i_4_ibuf (
    .O(desc_strproduct_addr_i_d[4]),
    .I(desc_strproduct_addr_i[4]) 
);
  IBUF desc_strproduct_addr_i_5_ibuf (
    .O(desc_strproduct_addr_i_d[5]),
    .I(desc_strproduct_addr_i[5]) 
);
  IBUF desc_strproduct_addr_i_6_ibuf (
    .O(desc_strproduct_addr_i_d[6]),
    .I(desc_strproduct_addr_i[6]) 
);
  IBUF desc_strproduct_addr_i_7_ibuf (
    .O(desc_strproduct_addr_i_d[7]),
    .I(desc_strproduct_addr_i[7]) 
);
  IBUF desc_strproduct_addr_i_8_ibuf (
    .O(desc_strproduct_addr_i_d[8]),
    .I(desc_strproduct_addr_i[8]) 
);
  IBUF desc_strproduct_addr_i_9_ibuf (
    .O(desc_strproduct_addr_i_d[9]),
    .I(desc_strproduct_addr_i[9]) 
);
  IBUF desc_strproduct_len_i_0_ibuf (
    .O(desc_strproduct_len_i_d[0]),
    .I(desc_strproduct_len_i[0]) 
);
  IBUF desc_strproduct_len_i_1_ibuf (
    .O(desc_strproduct_len_i_d[1]),
    .I(desc_strproduct_len_i[1]) 
);
  IBUF desc_strproduct_len_i_2_ibuf (
    .O(desc_strproduct_len_i_d[2]),
    .I(desc_strproduct_len_i[2]) 
);
  IBUF desc_strproduct_len_i_3_ibuf (
    .O(desc_strproduct_len_i_d[3]),
    .I(desc_strproduct_len_i[3]) 
);
  IBUF desc_strproduct_len_i_4_ibuf (
    .O(desc_strproduct_len_i_d[4]),
    .I(desc_strproduct_len_i[4]) 
);
  IBUF desc_strproduct_len_i_5_ibuf (
    .O(desc_strproduct_len_i_d[5]),
    .I(desc_strproduct_len_i[5]) 
);
  IBUF desc_strproduct_len_i_6_ibuf (
    .O(desc_strproduct_len_i_d[6]),
    .I(desc_strproduct_len_i[6]) 
);
  IBUF desc_strproduct_len_i_7_ibuf (
    .O(desc_strproduct_len_i_d[7]),
    .I(desc_strproduct_len_i[7]) 
);
  IBUF desc_strserial_addr_i_0_ibuf (
    .O(desc_strserial_addr_i_d[0]),
    .I(desc_strserial_addr_i[0]) 
);
  IBUF desc_strserial_addr_i_1_ibuf (
    .O(desc_strserial_addr_i_d[1]),
    .I(desc_strserial_addr_i[1]) 
);
  IBUF desc_strserial_addr_i_2_ibuf (
    .O(desc_strserial_addr_i_d[2]),
    .I(desc_strserial_addr_i[2]) 
);
  IBUF desc_strserial_addr_i_3_ibuf (
    .O(desc_strserial_addr_i_d[3]),
    .I(desc_strserial_addr_i[3]) 
);
  IBUF desc_strserial_addr_i_4_ibuf (
    .O(desc_strserial_addr_i_d[4]),
    .I(desc_strserial_addr_i[4]) 
);
  IBUF desc_strserial_addr_i_5_ibuf (
    .O(desc_strserial_addr_i_d[5]),
    .I(desc_strserial_addr_i[5]) 
);
  IBUF desc_strserial_addr_i_6_ibuf (
    .O(desc_strserial_addr_i_d[6]),
    .I(desc_strserial_addr_i[6]) 
);
  IBUF desc_strserial_addr_i_7_ibuf (
    .O(desc_strserial_addr_i_d[7]),
    .I(desc_strserial_addr_i[7]) 
);
  IBUF desc_strserial_addr_i_8_ibuf (
    .O(desc_strserial_addr_i_d[8]),
    .I(desc_strserial_addr_i[8]) 
);
  IBUF desc_strserial_addr_i_9_ibuf (
    .O(desc_strserial_addr_i_d[9]),
    .I(desc_strserial_addr_i[9]) 
);
  IBUF desc_strserial_len_i_0_ibuf (
    .O(desc_strserial_len_i_d[0]),
    .I(desc_strserial_len_i[0]) 
);
  IBUF desc_strserial_len_i_1_ibuf (
    .O(desc_strserial_len_i_d[1]),
    .I(desc_strserial_len_i[1]) 
);
  IBUF desc_strserial_len_i_2_ibuf (
    .O(desc_strserial_len_i_d[2]),
    .I(desc_strserial_len_i[2]) 
);
  IBUF desc_strserial_len_i_3_ibuf (
    .O(desc_strserial_len_i_d[3]),
    .I(desc_strserial_len_i[3]) 
);
  IBUF desc_strserial_len_i_4_ibuf (
    .O(desc_strserial_len_i_d[4]),
    .I(desc_strserial_len_i[4]) 
);
  IBUF desc_strserial_len_i_5_ibuf (
    .O(desc_strserial_len_i_d[5]),
    .I(desc_strserial_len_i[5]) 
);
  IBUF desc_strserial_len_i_6_ibuf (
    .O(desc_strserial_len_i_d[6]),
    .I(desc_strserial_len_i[6]) 
);
  IBUF desc_strserial_len_i_7_ibuf (
    .O(desc_strserial_len_i_d[7]),
    .I(desc_strserial_len_i[7]) 
);
  IBUF desc_have_strings_i_ibuf (
    .O(desc_have_strings_i_d),
    .I(desc_have_strings_i) 
);
  IBUF utmi_txready_i_ibuf (
    .O(utmi_txready_i_d),
    .I(utmi_txready_i) 
);
  IBUF utmi_datain_i_0_ibuf (
    .O(utmi_datain_i_d[0]),
    .I(utmi_datain_i[0]) 
);
  IBUF utmi_datain_i_1_ibuf (
    .O(utmi_datain_i_d[1]),
    .I(utmi_datain_i[1]) 
);
  IBUF utmi_datain_i_2_ibuf (
    .O(utmi_datain_i_d[2]),
    .I(utmi_datain_i[2]) 
);
  IBUF utmi_datain_i_3_ibuf (
    .O(utmi_datain_i_d[3]),
    .I(utmi_datain_i[3]) 
);
  IBUF utmi_datain_i_4_ibuf (
    .O(utmi_datain_i_d[4]),
    .I(utmi_datain_i[4]) 
);
  IBUF utmi_datain_i_5_ibuf (
    .O(utmi_datain_i_d[5]),
    .I(utmi_datain_i[5]) 
);
  IBUF utmi_datain_i_6_ibuf (
    .O(utmi_datain_i_d[6]),
    .I(utmi_datain_i[6]) 
);
  IBUF utmi_datain_i_7_ibuf (
    .O(utmi_datain_i_d[7]),
    .I(utmi_datain_i[7]) 
);
  IBUF utmi_rxactive_i_ibuf (
    .O(utmi_rxactive_i_d),
    .I(utmi_rxactive_i) 
);
  IBUF utmi_rxvalid_i_ibuf (
    .O(utmi_rxvalid_i_d),
    .I(utmi_rxvalid_i) 
);
  IBUF utmi_rxerror_i_ibuf (
    .O(utmi_rxerror_i_d),
    .I(utmi_rxerror_i) 
);
  IBUF utmi_linestate_i_0_ibuf (
    .O(utmi_linestate_i_d[0]),
    .I(utmi_linestate_i[0]) 
);
  IBUF utmi_linestate_i_1_ibuf (
    .O(utmi_linestate_i_d[1]),
    .I(utmi_linestate_i[1]) 
);
  OBUF usbrst_o_obuf (
    .O(usbrst_o),
    .I(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  OBUF highspeed_o_obuf (
    .O(highspeed_o),
    .I(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
  OBUF suspend_o_obuf (
    .O(suspend_o),
    .I(u_usb_device_controller_u_usb_init_suspend_o_d) 
);
  OBUF online_o_obuf (
    .O(online_o),
    .I(u_usb_device_controller_usb_control_inst_online_o_d) 
);
  OBUF txpop_o_obuf (
    .O(txpop_o),
    .I(u_usb_device_controller_usb_transact_inst_txpop_o_d) 
);
  OBUF txact_o_obuf (
    .O(txact_o),
    .I(u_usb_device_controller_txact_o_d) 
);
  OBUF txpktfin_o_obuf (
    .O(txpktfin_o),
    .I(u_usb_device_controller_txpktfin_o_d) 
);
  OBUF rxdat_o_0_obuf (
    .O(rxdat_o[0]),
    .I(u_usb_device_controller_rxdat_o_d[0]) 
);
  OBUF rxdat_o_1_obuf (
    .O(rxdat_o[1]),
    .I(u_usb_device_controller_rxdat_o_d[1]) 
);
  OBUF rxdat_o_2_obuf (
    .O(rxdat_o[2]),
    .I(u_usb_device_controller_rxdat_o_d[2]) 
);
  OBUF rxdat_o_3_obuf (
    .O(rxdat_o[3]),
    .I(u_usb_device_controller_rxdat_o_d[3]) 
);
  OBUF rxdat_o_4_obuf (
    .O(rxdat_o[4]),
    .I(u_usb_device_controller_rxdat_o_d[4]) 
);
  OBUF rxdat_o_5_obuf (
    .O(rxdat_o[5]),
    .I(u_usb_device_controller_rxdat_o_d[5]) 
);
  OBUF rxdat_o_6_obuf (
    .O(rxdat_o[6]),
    .I(u_usb_device_controller_rxdat_o_d[6]) 
);
  OBUF rxdat_o_7_obuf (
    .O(rxdat_o[7]),
    .I(u_usb_device_controller_rxdat_o_d[7]) 
);
  OBUF rxval_o_obuf (
    .O(rxval_o),
    .I(u_usb_device_controller_rxval_o_d) 
);
  OBUF rxact_o_obuf (
    .O(rxact_o),
    .I(u_usb_device_controller_rxact_o_d) 
);
  OBUF rxpktval_o_obuf (
    .O(rxpktval_o),
    .I(u_usb_device_controller_rxpktval_o_d) 
);
  OBUF setup_o_obuf (
    .O(setup_o),
    .I(u_usb_device_controller_setup_o_d) 
);
  OBUF endpt_o_0_obuf (
    .O(endpt_o[0]),
    .I(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
  OBUF endpt_o_1_obuf (
    .O(endpt_o[1]),
    .I(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  OBUF endpt_o_2_obuf (
    .O(endpt_o[2]),
    .I(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
  OBUF endpt_o_3_obuf (
    .O(endpt_o[3]),
    .I(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
  OBUF sof_o_obuf (
    .O(sof_o),
    .I(u_usb_device_controller_usb_transact_inst_sof_o_d) 
);
  OBUF inf_alter_o_0_obuf (
    .O(inf_alter_o[0]),
    .I(u_usb_device_controller_usb_control_inst_inf_alter_o_d[0]) 
);
  OBUF inf_alter_o_1_obuf (
    .O(inf_alter_o[1]),
    .I(u_usb_device_controller_usb_control_inst_inf_alter_o_d[1]) 
);
  OBUF inf_alter_o_2_obuf (
    .O(inf_alter_o[2]),
    .I(u_usb_device_controller_usb_control_inst_inf_alter_o_d[2]) 
);
  OBUF inf_alter_o_3_obuf (
    .O(inf_alter_o[3]),
    .I(u_usb_device_controller_usb_control_inst_inf_alter_o_d[3]) 
);
  OBUF inf_alter_o_4_obuf (
    .O(inf_alter_o[4]),
    .I(u_usb_device_controller_usb_control_inst_inf_alter_o_d[4]) 
);
  OBUF inf_alter_o_5_obuf (
    .O(inf_alter_o[5]),
    .I(u_usb_device_controller_usb_control_inst_inf_alter_o_d[5]) 
);
  OBUF inf_alter_o_6_obuf (
    .O(inf_alter_o[6]),
    .I(u_usb_device_controller_usb_control_inst_inf_alter_o_d[6]) 
);
  OBUF inf_alter_o_7_obuf (
    .O(inf_alter_o[7]),
    .I(u_usb_device_controller_usb_control_inst_inf_alter_o_d[7]) 
);
  OBUF inf_sel_o_0_obuf (
    .O(inf_sel_o[0]),
    .I(u_usb_device_controller_usb_control_inst_inf_sel_o_d[0]) 
);
  OBUF inf_sel_o_1_obuf (
    .O(inf_sel_o[1]),
    .I(u_usb_device_controller_usb_control_inst_inf_sel_o_d[1]) 
);
  OBUF inf_sel_o_2_obuf (
    .O(inf_sel_o[2]),
    .I(u_usb_device_controller_usb_control_inst_inf_sel_o_d[2]) 
);
  OBUF inf_sel_o_3_obuf (
    .O(inf_sel_o[3]),
    .I(u_usb_device_controller_usb_control_inst_inf_sel_o_d[3]) 
);
  OBUF inf_sel_o_4_obuf (
    .O(inf_sel_o[4]),
    .I(u_usb_device_controller_usb_control_inst_inf_sel_o_d[4]) 
);
  OBUF inf_sel_o_5_obuf (
    .O(inf_sel_o[5]),
    .I(u_usb_device_controller_usb_control_inst_inf_sel_o_d[5]) 
);
  OBUF inf_sel_o_6_obuf (
    .O(inf_sel_o[6]),
    .I(u_usb_device_controller_usb_control_inst_inf_sel_o_d[6]) 
);
  OBUF inf_sel_o_7_obuf (
    .O(inf_sel_o[7]),
    .I(u_usb_device_controller_usb_control_inst_inf_sel_o_d[7]) 
);
  OBUF inf_set_o_obuf (
    .O(inf_set_o),
    .I(u_usb_device_controller_usb_control_inst_inf_set_o_d) 
);
  OBUF descrom_raddr_o_0_obuf (
    .O(descrom_raddr_o[0]),
    .I(u_usb_device_controller_descrom_raddr_o_d[0]) 
);
  OBUF descrom_raddr_o_1_obuf (
    .O(descrom_raddr_o[1]),
    .I(u_usb_device_controller_descrom_raddr_o_d[1]) 
);
  OBUF descrom_raddr_o_2_obuf (
    .O(descrom_raddr_o[2]),
    .I(u_usb_device_controller_descrom_raddr_o_d[2]) 
);
  OBUF descrom_raddr_o_3_obuf (
    .O(descrom_raddr_o[3]),
    .I(u_usb_device_controller_descrom_raddr_o_d[3]) 
);
  OBUF descrom_raddr_o_4_obuf (
    .O(descrom_raddr_o[4]),
    .I(u_usb_device_controller_descrom_raddr_o_d[4]) 
);
  OBUF descrom_raddr_o_5_obuf (
    .O(descrom_raddr_o[5]),
    .I(u_usb_device_controller_descrom_raddr_o_d[5]) 
);
  OBUF descrom_raddr_o_6_obuf (
    .O(descrom_raddr_o[6]),
    .I(u_usb_device_controller_descrom_raddr_o_d[6]) 
);
  OBUF descrom_raddr_o_7_obuf (
    .O(descrom_raddr_o[7]),
    .I(u_usb_device_controller_descrom_raddr_o_d[7]) 
);
  OBUF descrom_raddr_o_8_obuf (
    .O(descrom_raddr_o[8]),
    .I(u_usb_device_controller_descrom_raddr_o_d[8]) 
);
  OBUF descrom_raddr_o_9_obuf (
    .O(descrom_raddr_o[9]),
    .I(u_usb_device_controller_descrom_raddr_o_d[9]) 
);
  OBUF utmi_dataout_o_0_obuf (
    .O(utmi_dataout_o[0]),
    .I(u_usb_device_controller_utmi_dataout_o_d[0]) 
);
  OBUF utmi_dataout_o_1_obuf (
    .O(utmi_dataout_o[1]),
    .I(u_usb_device_controller_utmi_dataout_o_d[1]) 
);
  OBUF utmi_dataout_o_2_obuf (
    .O(utmi_dataout_o[2]),
    .I(u_usb_device_controller_utmi_dataout_o_d[2]) 
);
  OBUF utmi_dataout_o_3_obuf (
    .O(utmi_dataout_o[3]),
    .I(u_usb_device_controller_utmi_dataout_o_d[3]) 
);
  OBUF utmi_dataout_o_4_obuf (
    .O(utmi_dataout_o[4]),
    .I(u_usb_device_controller_utmi_dataout_o_d[4]) 
);
  OBUF utmi_dataout_o_5_obuf (
    .O(utmi_dataout_o[5]),
    .I(u_usb_device_controller_utmi_dataout_o_d[5]) 
);
  OBUF utmi_dataout_o_6_obuf (
    .O(utmi_dataout_o[6]),
    .I(u_usb_device_controller_utmi_dataout_o_d[6]) 
);
  OBUF utmi_dataout_o_7_obuf (
    .O(utmi_dataout_o[7]),
    .I(u_usb_device_controller_utmi_dataout_o_d[7]) 
);
  OBUF utmi_txvalid_o_obuf (
    .O(utmi_txvalid_o),
    .I(u_usb_device_controller_utmi_txvalid_o_d) 
);
  OBUF utmi_opmode_o_0_obuf (
    .O(utmi_opmode_o[0]),
    .I(u_usb_device_controller_utmi_opmode_o_d[0]) 
);
  OBUF utmi_opmode_o_1_obuf (
    .O(utmi_opmode_o[1]),
    .I(u_usb_device_controller_utmi_opmode_o_d[1]) 
);
  OBUF utmi_xcvrselect_o_0_obuf (
    .O(utmi_xcvrselect_o[0]),
    .I(u_usb_device_controller_u_usb_init_utmi_xcvrselect_o_d[0]) 
);
  OBUF utmi_xcvrselect_o_1_obuf (
    .O(utmi_xcvrselect_o[1]),
    .I(GND) 
);
  OBUF utmi_termselect_o_obuf (
    .O(utmi_termselect_o),
    .I(u_usb_device_controller_u_usb_init_utmi_termselect_o_d) 
);
  OBUF utmi_reset_o_obuf (
    .O(utmi_reset_o),
    .I(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFR \u_usb_device_controller/s_endpt_rxrdy_s0  (
    .Q(u_usb_device_controller_s_endpt_rxrdy),
    .D(rxrdy_i_d),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/s_endpt_txcork_s0  (
    .Q(u_usb_device_controller_s_endpt_txcork),
    .D(u_usb_device_controller_n1240),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/s_halt_out_s0  (
    .Q(u_usb_device_controller_s_halt_out),
    .D(u_usb_device_controller_n1241),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/s_halt_in_s0  (
    .Q(u_usb_device_controller_s_halt_in),
    .D(u_usb_device_controller_n1242),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/s_osync_s0  (
    .Q(u_usb_device_controller_s_osync),
    .D(u_usb_device_controller_n1243),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/s_isync_s0  (
    .Q(u_usb_device_controller_s_isync),
    .D(u_usb_device_controller_n1244),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_11_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[11]),
    .D(txdat_len_i_d[11]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_10_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[10]),
    .D(u_usb_device_controller_n1261),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_9_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[9]),
    .D(txdat_len_i_d[9]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_8_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[8]),
    .D(txdat_len_i_d[8]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_7_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[7]),
    .D(txdat_len_i_d[7]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_6_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[6]),
    .D(txdat_len_i_d[6]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFS \u_usb_device_controller/s_txbuf_stop_5_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[5]),
    .D(u_usb_device_controller_n1266),
    .CLK(clk_i_d),
    .SET(reset_i_d) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_4_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[4]),
    .D(txdat_len_i_d[4]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_3_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[3]),
    .D(txdat_len_i_d[3]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_2_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[2]),
    .D(txdat_len_i_d[2]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_1_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[1]),
    .D(txdat_len_i_d[1]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFR \u_usb_device_controller/s_txbuf_stop_0_s0  (
    .Q(u_usb_device_controller_s_txbuf_stop[0]),
    .D(txdat_len_i_d[0]),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2339) 
);
  DFFR \u_usb_device_controller/cur_state_3_s0  (
    .Q(u_usb_device_controller_cur_state[3]),
    .D(u_usb_device_controller_next_state[3]),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/cur_state_2_s0  (
    .Q(u_usb_device_controller_cur_state[2]),
    .D(u_usb_device_controller_next_state[2]),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/cur_state_1_s0  (
    .Q(u_usb_device_controller_cur_state[1]),
    .D(u_usb_device_controller_next_state[1]),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFR \u_usb_device_controller/cur_state_0_s0  (
    .Q(u_usb_device_controller_cur_state[0]),
    .D(u_usb_device_controller_next_state[0]),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
  DFFC \u_usb_device_controller/rxdat_d2_7_s0  (
    .Q(u_usb_device_controller_rxdat_d2[7]),
    .D(u_usb_device_controller_n1760),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFC \u_usb_device_controller/rxdat_d2_6_s0  (
    .Q(u_usb_device_controller_rxdat_d2[6]),
    .D(u_usb_device_controller_n1761),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFC \u_usb_device_controller/rxdat_d2_5_s0  (
    .Q(u_usb_device_controller_rxdat_d2[5]),
    .D(u_usb_device_controller_n1762),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFC \u_usb_device_controller/rxdat_d2_4_s0  (
    .Q(u_usb_device_controller_rxdat_d2[4]),
    .D(u_usb_device_controller_n1763),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFC \u_usb_device_controller/rxdat_d2_3_s0  (
    .Q(u_usb_device_controller_rxdat_d2[3]),
    .D(u_usb_device_controller_n1764),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFC \u_usb_device_controller/rxdat_d2_2_s0  (
    .Q(u_usb_device_controller_rxdat_d2[2]),
    .D(u_usb_device_controller_n1765),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFC \u_usb_device_controller/rxdat_d2_1_s0  (
    .Q(u_usb_device_controller_rxdat_d2[1]),
    .D(u_usb_device_controller_n1766),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFC \u_usb_device_controller/rxdat_d2_0_s0  (
    .Q(u_usb_device_controller_rxdat_d2[0]),
    .D(u_usb_device_controller_n1767),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFC \u_usb_device_controller/rxval_d2_s0  (
    .Q(u_usb_device_controller_rxval_d2),
    .D(u_usb_device_controller_n1770),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFC \u_usb_device_controller/rx_packet_valid_s0  (
    .Q(u_usb_device_controller_rxpktval_o_d),
    .D(u_usb_device_controller_n1810),
    .CLK(clk_i_d),
    .CLEAR(reset_i_d) 
);
  DFFE \u_usb_device_controller/descrom_raddr_9_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[9]),
    .D(u_usb_device_controller_n2024),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFE \u_usb_device_controller/descrom_raddr_8_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[8]),
    .D(u_usb_device_controller_n2025),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFE \u_usb_device_controller/descrom_raddr_7_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[7]),
    .D(u_usb_device_controller_n2026),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFE \u_usb_device_controller/descrom_raddr_6_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[6]),
    .D(u_usb_device_controller_n2027),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFE \u_usb_device_controller/descrom_raddr_5_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[5]),
    .D(u_usb_device_controller_n2028),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFE \u_usb_device_controller/descrom_raddr_4_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[4]),
    .D(u_usb_device_controller_n2029),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFE \u_usb_device_controller/descrom_raddr_3_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[3]),
    .D(u_usb_device_controller_n2030),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFE \u_usb_device_controller/descrom_raddr_2_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[2]),
    .D(u_usb_device_controller_n2031),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFE \u_usb_device_controller/descrom_raddr_1_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[1]),
    .D(u_usb_device_controller_n2032),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFE \u_usb_device_controller/descrom_raddr_0_s0  (
    .Q(u_usb_device_controller_descrom_raddr_o_d[0]),
    .D(u_usb_device_controller_n2033),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_dscrd) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_en_dly_s0  (
    .Q(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .D(VCC),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_n378),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_en_dect_s0  (
    .Q(u_usb_device_controller_test_packet_inst_test_en_dect),
    .D(VCC),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_usbc_test_en),
    .CLEAR(reset_i_d) 
);
  DFFS \u_usb_device_controller/u_usb_init/v_clrtimer2_s0  (
    .Q(u_usb_device_controller_u_usb_init_v_clrtimer2),
    .D(u_usb_device_controller_u_usb_init_n212),
    .CLK(clk_i_d),
    .SET(reset_i_d) 
);
  DFF \u_usb_device_controller/u_usb_init/s_linestate_1_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_linestate[1]),
    .D(utmi_linestate_i_d[1]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_init/s_linestate_0_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .D(utmi_linestate_i_d[0]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_init/s_usb_test_en_0_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_usb_test_en[0]),
    .D(u_usb_device_controller_usb_control_inst_usbc_test_en),
    .CLK(clk_i_d) 
);
  DFFS \u_usb_device_controller/u_usb_init/s_reset_s0  (
    .Q(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .D(u_usb_device_controller_u_usb_init_n213),
    .CLK(clk_i_d),
    .SET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_reset_s0 .INIT=1'b1;
  DFFR \u_usb_device_controller/u_usb_init/s_chirpk_s0  (
    .Q(u_usb_device_controller_u_usb_init_usbp_chirpk),
    .D(u_usb_device_controller_u_usb_init_n223),
    .CLK(clk_i_d),
    .RESET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpk_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_highspeed_s0  (
    .Q(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .D(u_usb_device_controller_u_usb_init_n218),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_highspeed),
    .RESET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_highspeed_s0 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_chirpcnt[2]),
    .D(u_usb_device_controller_u_usb_init_n220),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_chirpcnt_2) 
);
  DFFE \u_usb_device_controller/u_usb_init/s_chirpcnt_1_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_chirpcnt[1]),
    .D(u_usb_device_controller_u_usb_init_n221),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_chirpcnt_2) 
);
  DFFE \u_usb_device_controller/u_usb_init/s_chirpcnt_0_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_chirpcnt[0]),
    .D(u_usb_device_controller_u_usb_init_n222),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_chirpcnt_2) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_15_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[15]),
    .D(u_usb_device_controller_u_usb_init_n226),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_14_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[14]),
    .D(u_usb_device_controller_u_usb_init_n227),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_13_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[13]),
    .D(u_usb_device_controller_u_usb_init_n228),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_12_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[12]),
    .D(u_usb_device_controller_u_usb_init_n229),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_11_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[11]),
    .D(u_usb_device_controller_u_usb_init_n230),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_10_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[10]),
    .D(u_usb_device_controller_u_usb_init_n231),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_9_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[9]),
    .D(u_usb_device_controller_u_usb_init_n232),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_8_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[8]),
    .D(u_usb_device_controller_u_usb_init_n233),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_7_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[7]),
    .D(u_usb_device_controller_u_usb_init_n234),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_6_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[6]),
    .D(u_usb_device_controller_u_usb_init_n235),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_5_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[5]),
    .D(u_usb_device_controller_u_usb_init_n236),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_4_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[4]),
    .D(u_usb_device_controller_u_usb_init_n237),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_3_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[3]),
    .D(u_usb_device_controller_u_usb_init_n238),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_2_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[2]),
    .D(u_usb_device_controller_u_usb_init_n239),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer1_1_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[1]),
    .D(u_usb_device_controller_u_usb_init_n240),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_19_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[19]),
    .D(u_usb_device_controller_u_usb_init_n260),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_19_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_18_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[18]),
    .D(u_usb_device_controller_u_usb_init_n261),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_18_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_17_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[17]),
    .D(u_usb_device_controller_u_usb_init_n262),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_17_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_16_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[16]),
    .D(u_usb_device_controller_u_usb_init_n263),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_16_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_15_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[15]),
    .D(u_usb_device_controller_u_usb_init_n264),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_15_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_14_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[14]),
    .D(u_usb_device_controller_u_usb_init_n265),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_14_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_13_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[13]),
    .D(u_usb_device_controller_u_usb_init_n266),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_13_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_12_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[12]),
    .D(u_usb_device_controller_u_usb_init_n267),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_12_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_11_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[11]),
    .D(u_usb_device_controller_u_usb_init_n268),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_11_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_10_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[10]),
    .D(u_usb_device_controller_u_usb_init_n269),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_10_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_9_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[9]),
    .D(u_usb_device_controller_u_usb_init_n270),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_9_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_8_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[8]),
    .D(u_usb_device_controller_u_usb_init_n271),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_8_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_7_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[7]),
    .D(u_usb_device_controller_u_usb_init_n272),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_7_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_6_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[6]),
    .D(u_usb_device_controller_u_usb_init_n273),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_6_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_5_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[5]),
    .D(u_usb_device_controller_u_usb_init_n274),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_5_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_4_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[4]),
    .D(u_usb_device_controller_u_usb_init_n275),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_4_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_3_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[3]),
    .D(u_usb_device_controller_u_usb_init_n276),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_3_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_2_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[2]),
    .D(u_usb_device_controller_u_usb_init_n277),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_2_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_timer2_1_s0  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[1]),
    .D(u_usb_device_controller_u_usb_init_n278),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n316),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_1_s0 .INIT=1'b0;
  DFFCE \u_usb_device_controller/u_usb_init/s_suspend_s0  (
    .Q(u_usb_device_controller_u_usb_init_suspend_o_d),
    .D(VCC),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_n414),
    .CLEAR(u_usb_device_controller_u_usb_init_phy_linestate_rst) 
);
defparam \u_usb_device_controller/u_usb_init/s_suspend_s0 .INIT=1'b0;
  DFFS \u_usb_device_controller/u_usb_init/v_clrtimer1_s0  (
    .Q(u_usb_device_controller_u_usb_init_v_clrtimer1),
    .D(u_usb_device_controller_u_usb_init_n219),
    .CLK(clk_i_d),
    .SET(reset_i_d) 
);
  DFFR \u_usb_device_controller/u_usb_packet/s_txfirst_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_txfirst),
    .D(u_usb_device_controller_u_usb_packet_n328),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_u_usb_packet_n800) 
);
defparam \u_usb_device_controller/u_usb_packet/s_txfirst_s0 .INIT=1'b0;
  DFF \u_usb_device_controller/u_usb_packet/s_rxactive_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .D(utmi_rxactive_i_d),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_rxvalid_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .D(utmi_rxvalid_i_d),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_rxerror_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_rxerror),
    .D(utmi_rxerror_i_d),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_datain_7_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .D(utmi_datain_i_d[7]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_datain_6_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]),
    .D(utmi_datain_i_d[6]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_datain_5_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .D(utmi_datain_i_d[5]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_datain_4_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .D(utmi_datain_i_d[4]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_datain_3_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .D(utmi_datain_i_d[3]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_datain_2_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .D(utmi_datain_i_d[2]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_datain_1_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .D(utmi_datain_i_d[1]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_datain_0_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .D(utmi_datain_i_d[0]),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_txready_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_txready),
    .D(utmi_txready_i_d),
    .CLK(clk_i_d) 
);
  DFF \u_usb_device_controller/u_usb_packet/s_rxgoodpacket_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_rxgoodpacket),
    .D(u_usb_device_controller_u_usb_packet_n912),
    .CLK(clk_i_d) 
);
  DFFE \u_usb_device_controller/u_usb_packet/crc5_buf_4_s0  (
    .Q(u_usb_device_controller_u_usb_packet_crc5_buf[4]),
    .D(u_usb_device_controller_u_usb_packet_n571),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc5_buf_4) 
);
  DFFE \u_usb_device_controller/u_usb_packet/crc5_buf_3_s0  (
    .Q(u_usb_device_controller_u_usb_packet_crc5_buf[3]),
    .D(u_usb_device_controller_u_usb_packet_n573),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc5_buf_4) 
);
  DFFE \u_usb_device_controller/u_usb_packet/crc5_buf_2_s0  (
    .Q(u_usb_device_controller_u_usb_packet_crc5_buf[2]),
    .D(u_usb_device_controller_u_usb_packet_n575),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc5_buf_4) 
);
  DFFE \u_usb_device_controller/u_usb_packet/crc5_buf_1_s0  (
    .Q(u_usb_device_controller_u_usb_packet_crc5_buf[1]),
    .D(u_usb_device_controller_u_usb_packet_n577),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc5_buf_4) 
);
  DFFE \u_usb_device_controller/u_usb_packet/crc5_buf_0_s0  (
    .Q(u_usb_device_controller_u_usb_packet_crc5_buf[0]),
    .D(u_usb_device_controller_u_usb_packet_n579),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc5_buf_4) 
);
  DFFRE \u_usb_device_controller/u_usb_packet/PHY_DATAOUT_7_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_dataout_o[7]),
    .D(u_usb_device_controller_u_usb_packet_n778),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n919),
    .RESET(u_usb_device_controller_u_usb_packet_n1454) 
);
  DFFRE \u_usb_device_controller/u_usb_packet/PHY_DATAOUT_6_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_dataout_o[6]),
    .D(u_usb_device_controller_u_usb_packet_n779),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n919),
    .RESET(u_usb_device_controller_u_usb_packet_n1454) 
);
  DFFRE \u_usb_device_controller/u_usb_packet/PHY_DATAOUT_5_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_dataout_o[5]),
    .D(u_usb_device_controller_u_usb_packet_n780),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n919),
    .RESET(u_usb_device_controller_u_usb_packet_n1454) 
);
  DFFRE \u_usb_device_controller/u_usb_packet/PHY_DATAOUT_4_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_dataout_o[4]),
    .D(u_usb_device_controller_u_usb_packet_n781),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n919),
    .RESET(u_usb_device_controller_u_usb_packet_n1454) 
);
  DFFRE \u_usb_device_controller/u_usb_packet/PHY_DATAOUT_3_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_dataout_o[3]),
    .D(u_usb_device_controller_u_usb_packet_n782),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n919),
    .RESET(u_usb_device_controller_u_usb_packet_n1454) 
);
  DFFRE \u_usb_device_controller/u_usb_packet/PHY_DATAOUT_2_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_dataout_o[2]),
    .D(u_usb_device_controller_u_usb_packet_n783),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n919),
    .RESET(u_usb_device_controller_u_usb_packet_n1454) 
);
  DFFRE \u_usb_device_controller/u_usb_packet/PHY_DATAOUT_1_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_dataout_o[1]),
    .D(u_usb_device_controller_u_usb_packet_n784),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n919),
    .RESET(u_usb_device_controller_u_usb_packet_n1454) 
);
  DFFRE \u_usb_device_controller/u_usb_packet/PHY_DATAOUT_0_s0  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_dataout_o[0]),
    .D(u_usb_device_controller_u_usb_packet_n785),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n919),
    .RESET(u_usb_device_controller_u_usb_packet_n1454) 
);
  DFFE \u_usb_device_controller/u_usb_packet/s_dataout_7_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_dataout[7]),
    .D(u_usb_device_controller_u_usb_packet_n640),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
  DFFE \u_usb_device_controller/u_usb_packet/s_dataout_6_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_dataout[6]),
    .D(u_usb_device_controller_u_usb_packet_n642),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
  DFFE \u_usb_device_controller/u_usb_packet/s_dataout_5_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_dataout[5]),
    .D(u_usb_device_controller_u_usb_packet_n644),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
  DFFE \u_usb_device_controller/u_usb_packet/s_dataout_4_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_dataout[4]),
    .D(u_usb_device_controller_u_usb_packet_n646),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
  DFFE \u_usb_device_controller/u_usb_packet/s_dataout_3_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_dataout[3]),
    .D(u_usb_device_controller_u_usb_packet_n648),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
  DFFE \u_usb_device_controller/u_usb_packet/s_dataout_2_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_dataout[2]),
    .D(u_usb_device_controller_u_usb_packet_n650),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
  DFFE \u_usb_device_controller/u_usb_packet/s_dataout_1_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_dataout[1]),
    .D(u_usb_device_controller_u_usb_packet_n652),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
  DFFE \u_usb_device_controller/u_usb_packet/s_dataout_0_s0  (
    .Q(u_usb_device_controller_u_usb_packet_s_dataout[0]),
    .D(u_usb_device_controller_u_usb_packet_n654),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
  DFFR \u_usb_device_controller/usb_transact_inst/s_setup_s1  (
    .Q(u_usb_device_controller_usb_transact_inst_s_setup),
    .D(u_usb_device_controller_usb_transact_inst_n1068),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_transact_inst/s_endpt_3_s0  (
    .Q(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_s_endpt_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_endpt_3_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_endpt_2_s0  (
    .Q(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_s_endpt_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_endpt_2_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_endpt_1_s0  (
    .Q(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_s_endpt_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_endpt_1_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_endpt_0_s0  (
    .Q(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_s_endpt_0),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_endpt_0_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_osync_s0  (
    .Q(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1565),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_osync_s0 .INIT=1'b0;
  DFF \u_usb_device_controller/usb_transact_inst/s_prevrxact_s0  (
    .Q(u_usb_device_controller_usb_transact_inst_s_prevrxact),
    .D(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .CLK(clk_i_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_addr_6_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_addr[6]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[6]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2896),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_addr_6_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_addr_5_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_addr[5]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[5]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2896),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_addr_5_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_addr_4_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_addr[4]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[4]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2896),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_addr_4_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_addr_3_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_addr[3]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2896),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_addr_3_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_addr_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_addr[2]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2896),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_addr_2_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_addr_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_addr[1]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2896),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_addr_1_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_addr_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_addr[0]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2896),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_addr_0_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_confd_s0  (
    .Q(u_usb_device_controller_usb_control_inst_online_o_d),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1876),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_confd_s0 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_testmode_7_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_testmode[7]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1909),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_testmode_6_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_testmode[6]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[6]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1909),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_testmode_5_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_testmode[5]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[5]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1909),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_testmode_4_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_testmode[4]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[4]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1909),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_testmode_3_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_testmode[3]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1909),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_testmode_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_testmode[2]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1909),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_testmode_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_testmode[1]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1909),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_testmode_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .D(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1909),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_test_en_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_test_en),
    .D(VCC),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2902),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_test_sel_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_test_sel),
    .D(VCC),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1836),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_alter_7_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_alter_o_d[7]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1864),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_alter_6_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_alter_o_d[6]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1864),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_alter_5_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_alter_o_d[5]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1864),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_alter_4_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_alter_o_d[4]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1864),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_alter_3_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_alter_o_d[3]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1864),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_alter_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_alter_o_d[2]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1864),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_alter_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_alter_o_d[1]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1864),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_alter_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_alter_o_d[0]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1864),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_7_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_sel_o_d[7]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1837),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_6_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_sel_o_d[6]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1837),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_5_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_sel_o_d[5]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1837),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_4_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_sel_o_d[4]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1837),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_3_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_sel_o_d[3]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1837),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_sel_o_d[2]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1837),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_sel_o_d[1]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1837),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_inf_sel_o_d[0]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1837),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerptr_7_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscoff[7]),
    .D(u_usb_device_controller_usb_control_inst_n1617),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerptr_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerptr_6_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscoff[6]),
    .D(u_usb_device_controller_usb_control_inst_n1646),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerptr_7_8) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerptr_5_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscoff[5]),
    .D(u_usb_device_controller_usb_control_inst_n1649),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerptr_5) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerptr_4_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscoff[4]),
    .D(u_usb_device_controller_usb_control_inst_n1652),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerptr_5) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerptr_3_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscoff[3]),
    .D(u_usb_device_controller_usb_control_inst_n1655),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerptr_5) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerptr_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscoff[2]),
    .D(u_usb_device_controller_usb_control_inst_n1658),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerptr_5) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerptr_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]),
    .D(u_usb_device_controller_usb_control_inst_n1661),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerptr_5) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerptr_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .D(u_usb_device_controller_usb_control_inst_n1664),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerptr_5) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_setupptr_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .D(u_usb_device_controller_usb_control_inst_n1693),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_setupptr_2) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_setupptr_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .D(u_usb_device_controller_usb_control_inst_n1696),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_setupptr_2) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerlen_7_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_answerlen[7]),
    .D(u_usb_device_controller_usb_control_inst_n407),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerlen_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerlen_6_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_answerlen[6]),
    .D(u_usb_device_controller_usb_control_inst_n408),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerlen_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerlen_5_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_answerlen[5]),
    .D(u_usb_device_controller_usb_control_inst_n409),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerlen_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerlen_4_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_answerlen[4]),
    .D(u_usb_device_controller_usb_control_inst_n410),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerlen_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerlen_3_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_answerlen[3]),
    .D(u_usb_device_controller_usb_control_inst_n411),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerlen_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerlen_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_answerlen[2]),
    .D(u_usb_device_controller_usb_control_inst_n412),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerlen_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerlen_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_answerlen[1]),
    .D(u_usb_device_controller_usb_control_inst_n413),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerlen_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_answerlen_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_answerlen[0]),
    .D(u_usb_device_controller_usb_control_inst_n414),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_answerlen_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlparam_7_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .D(u_usb_device_controller_usb_control_inst_n435),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_ctlparam_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlparam_6_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscinx[6]),
    .D(u_usb_device_controller_usb_control_inst_n436),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_ctlparam_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlparam_5_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscinx[5]),
    .D(u_usb_device_controller_usb_control_inst_n437),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_ctlparam_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlparam_4_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscinx[4]),
    .D(u_usb_device_controller_usb_control_inst_n438),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_ctlparam_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlparam_3_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .D(u_usb_device_controller_usb_control_inst_n439),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_ctlparam_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlparam_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .D(u_usb_device_controller_usb_control_inst_n440),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_ctlparam_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlparam_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .D(u_usb_device_controller_usb_control_inst_n441),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_ctlparam_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlparam_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .D(u_usb_device_controller_usb_control_inst_n442),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_ctlparam_7) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_txdat[7]),
    .D(u_usb_device_controller_usb_control_inst_n1382),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_sendbyte_1) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s0 .INIT=1'b0;
  DFFE \u_usb_device_controller/usb_control_inst/s_sendbyte_6_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_txdat[6]),
    .D(u_usb_device_controller_usb_control_inst_n1383),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_sendbyte_1) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_6_s0 .INIT=1'b0;
  DFFE \u_usb_device_controller/usb_control_inst/s_sendbyte_5_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_txdat[5]),
    .D(u_usb_device_controller_usb_control_inst_n1384),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_sendbyte_1) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_5_s0 .INIT=1'b0;
  DFFE \u_usb_device_controller/usb_control_inst/s_sendbyte_4_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_txdat[4]),
    .D(u_usb_device_controller_usb_control_inst_n1385),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_sendbyte_1) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_4_s0 .INIT=1'b0;
  DFFE \u_usb_device_controller/usb_control_inst/s_sendbyte_3_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_txdat[3]),
    .D(u_usb_device_controller_usb_control_inst_n1386),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_sendbyte_1) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_3_s0 .INIT=1'b0;
  DFFE \u_usb_device_controller/usb_control_inst/s_sendbyte_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_txdat[2]),
    .D(u_usb_device_controller_usb_control_inst_n1387),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_sendbyte_1) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_2_s0 .INIT=1'b0;
  DFFE \u_usb_device_controller/usb_control_inst/s_sendbyte_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_txdat[1]),
    .D(u_usb_device_controller_usb_control_inst_n1388),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_sendbyte_1) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_1_s0 .INIT=1'b0;
  DFFE \u_usb_device_controller/usb_control_inst/s_sendbyte_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_txdat[0]),
    .D(u_usb_device_controller_usb_control_inst_n1860),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_sendbyte_7) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_0_s0 .INIT=1'b0;
  DFFE \u_usb_device_controller/usb_control_inst/s_desctyp_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2067) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_desctyp_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2067) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_desctyp_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2067) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlrequest_3_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2070) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlrequest_2_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2070) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlrequest_1_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2070) 
);
  DFFE \u_usb_device_controller/usb_control_inst/s_ctlrequest_0_s0  (
    .Q(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .D(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n2070) 
);
  DLC \u_usb_device_controller/next_state_3_s0  (
    .Q(u_usb_device_controller_next_state[3]),
    .D(u_usb_device_controller_n1519),
    .G(u_usb_device_controller_n1520),
    .CLEAR(u_usb_device_controller_n2219) 
);
  DLC \u_usb_device_controller/next_state_2_s0  (
    .Q(u_usb_device_controller_next_state[2]),
    .D(u_usb_device_controller_n1524),
    .G(u_usb_device_controller_n1520),
    .CLEAR(u_usb_device_controller_n2219) 
);
  DLC \u_usb_device_controller/next_state_1_s0  (
    .Q(u_usb_device_controller_next_state[1]),
    .D(u_usb_device_controller_n1529),
    .G(u_usb_device_controller_n1520),
    .CLEAR(u_usb_device_controller_n2219) 
);
  DLC \u_usb_device_controller/next_state_0_s0  (
    .Q(u_usb_device_controller_next_state[0]),
    .D(u_usb_device_controller_n1534),
    .G(u_usb_device_controller_n1520),
    .CLEAR(u_usb_device_controller_n2219) 
);
  DFFCE \u_usb_device_controller/rxdat_d0_7_s1  (
    .Q(u_usb_device_controller_rxdat_d0[7]),
    .D(u_usb_device_controller_n1699),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d0_7_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d0_6_s1  (
    .Q(u_usb_device_controller_rxdat_d0[6]),
    .D(u_usb_device_controller_n1700),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d0_6_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d0_5_s1  (
    .Q(u_usb_device_controller_rxdat_d0[5]),
    .D(u_usb_device_controller_n1701),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d0_5_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d0_4_s1  (
    .Q(u_usb_device_controller_rxdat_d0[4]),
    .D(u_usb_device_controller_n1702),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d0_4_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d0_3_s1  (
    .Q(u_usb_device_controller_rxdat_d0[3]),
    .D(u_usb_device_controller_n1703),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d0_3_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d0_2_s1  (
    .Q(u_usb_device_controller_rxdat_d0[2]),
    .D(u_usb_device_controller_n1704),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d0_2_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d0_1_s1  (
    .Q(u_usb_device_controller_rxdat_d0[1]),
    .D(u_usb_device_controller_n1705),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d0_1_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d0_0_s1  (
    .Q(u_usb_device_controller_rxdat_d0[0]),
    .D(u_usb_device_controller_n1706),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d0_0_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d1_7_s1  (
    .Q(u_usb_device_controller_rxdat_d1[7]),
    .D(u_usb_device_controller_n1707),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d1_7_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d1_6_s1  (
    .Q(u_usb_device_controller_rxdat_d1[6]),
    .D(u_usb_device_controller_n1708),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d1_6_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d1_5_s1  (
    .Q(u_usb_device_controller_rxdat_d1[5]),
    .D(u_usb_device_controller_n1709),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d1_5_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d1_4_s1  (
    .Q(u_usb_device_controller_rxdat_d1[4]),
    .D(u_usb_device_controller_n1710),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d1_4_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d1_3_s1  (
    .Q(u_usb_device_controller_rxdat_d1[3]),
    .D(u_usb_device_controller_n1711),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d1_3_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d1_2_s1  (
    .Q(u_usb_device_controller_rxdat_d1[2]),
    .D(u_usb_device_controller_n1712),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d1_2_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d1_1_s1  (
    .Q(u_usb_device_controller_rxdat_d1[1]),
    .D(u_usb_device_controller_n1713),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d1_1_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxdat_d1_0_s1  (
    .Q(u_usb_device_controller_rxdat_d1[0]),
    .D(u_usb_device_controller_n1714),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxdat_d1_0_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxval_d0_s1  (
    .Q(u_usb_device_controller_rxval_d0),
    .D(u_usb_device_controller_n2393),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxval_d0_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/rxval_d1_s1  (
    .Q(u_usb_device_controller_rxval_d1),
    .D(u_usb_device_controller_n1716),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_rxdat_d0_7),
    .CLEAR(reset_i_d) 
);
defparam \u_usb_device_controller/rxval_d1_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_opmode_1_s1  (
    .Q(u_usb_device_controller_u_usb_init_usbi_opmode[1]),
    .D(u_usb_device_controller_u_usb_init_n208),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_opmode_0),
    .RESET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_opmode_1_s1 .INIT=1'b0;
  DFFSE \u_usb_device_controller/u_usb_init/s_opmode_0_s1  (
    .Q(u_usb_device_controller_u_usb_init_usbi_opmode[0]),
    .D(u_usb_device_controller_u_usb_init_n209),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_opmode_0),
    .SET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_opmode_0_s1 .INIT=1'b1;
  DFFSE \u_usb_device_controller/u_usb_init/s_xcvrselect_s1  (
    .Q(u_usb_device_controller_u_usb_init_utmi_xcvrselect_o_d[0]),
    .D(u_usb_device_controller_u_usb_init_n210),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_opmode_0),
    .SET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_xcvrselect_s1 .INIT=1'b1;
  DFFSE \u_usb_device_controller/u_usb_init/s_termselect_s1  (
    .Q(u_usb_device_controller_u_usb_init_utmi_termselect_o_d),
    .D(u_usb_device_controller_u_usb_init_n211),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_opmode_0),
    .SET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_termselect_s1 .INIT=1'b1;
  DFFRE \u_usb_device_controller/u_usb_init/s_state_3_s1  (
    .Q(u_usb_device_controller_u_usb_init_s_state[3]),
    .D(u_usb_device_controller_u_usb_init_n214),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_state_0),
    .RESET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_15_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[15]),
    .D(u_usb_device_controller_u_usb_packet_n761),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_15_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_14_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[14]),
    .D(u_usb_device_controller_u_usb_packet_n762),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_14_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_13_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[13]),
    .D(u_usb_device_controller_u_usb_packet_n763),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_13_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_12_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[12]),
    .D(u_usb_device_controller_u_usb_packet_n764),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_12_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_11_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[11]),
    .D(u_usb_device_controller_u_usb_packet_n765),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_11_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_10_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[10]),
    .D(u_usb_device_controller_u_usb_packet_n766),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_10_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_9_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[9]),
    .D(u_usb_device_controller_u_usb_packet_n767),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_9_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_8_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[8]),
    .D(u_usb_device_controller_u_usb_packet_n768),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_8_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_7_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[7]),
    .D(u_usb_device_controller_u_usb_packet_n769),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_7_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_6_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[6]),
    .D(u_usb_device_controller_u_usb_packet_n770),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_6_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_5_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[5]),
    .D(u_usb_device_controller_u_usb_packet_n771),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_5_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_4_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[4]),
    .D(u_usb_device_controller_u_usb_packet_n772),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_4_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_3_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[3]),
    .D(u_usb_device_controller_u_usb_packet_n773),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_3_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_2_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[2]),
    .D(u_usb_device_controller_u_usb_packet_n774),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_2_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_1_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[1]),
    .D(u_usb_device_controller_u_usb_packet_n775),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_1_s1 .INIT=1'b0;
  DFFE \u_usb_device_controller/u_usb_packet/crc16_buf_0_s1  (
    .Q(u_usb_device_controller_u_usb_packet_crc16_buf[0]),
    .D(u_usb_device_controller_u_usb_packet_n776),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_crc16_buf_15) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_0_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/PHY_TXVALID_s1  (
    .Q(u_usb_device_controller_u_usb_packet_usbp_txvalid_o),
    .D(u_usb_device_controller_u_usb_packet_n920),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_PHY_TXVALID),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/PHY_TXVALID_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_11_s2  (
    .Q(u_usb_device_controller_s_bufptr[11]),
    .D(u_usb_device_controller_n1593),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_11_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_10_s2  (
    .Q(u_usb_device_controller_s_bufptr[10]),
    .D(u_usb_device_controller_n1595),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_10_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_9_s2  (
    .Q(u_usb_device_controller_s_bufptr[9]),
    .D(u_usb_device_controller_n1597),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_9_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_8_s2  (
    .Q(u_usb_device_controller_s_bufptr[8]),
    .D(u_usb_device_controller_n1599),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_8_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_7_s2  (
    .Q(u_usb_device_controller_s_bufptr[7]),
    .D(u_usb_device_controller_n1601),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_7_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_6_s2  (
    .Q(u_usb_device_controller_s_bufptr[6]),
    .D(u_usb_device_controller_n1603),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_6_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_5_s2  (
    .Q(u_usb_device_controller_s_bufptr[5]),
    .D(u_usb_device_controller_n1605),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_5_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_4_s2  (
    .Q(u_usb_device_controller_s_bufptr[4]),
    .D(u_usb_device_controller_n1607),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_4_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_3_s2  (
    .Q(u_usb_device_controller_s_bufptr[3]),
    .D(u_usb_device_controller_n1609),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_3_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_2_s2  (
    .Q(u_usb_device_controller_s_bufptr[2]),
    .D(u_usb_device_controller_n1611),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_2_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_1_s2  (
    .Q(u_usb_device_controller_s_bufptr[1]),
    .D(u_usb_device_controller_n1613),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_bufptr_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_1_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_bufptr_0_s2  (
    .Q(u_usb_device_controller_s_bufptr[0]),
    .D(u_usb_device_controller_n1615),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n1593_24),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_bufptr_0_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_endpt_tx_en_s1  (
    .Q(u_usb_device_controller_txact_o_d),
    .D(u_usb_device_controller_n1585),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n1619),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_endpt_tx_en_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/s_nyet_s2  (
    .Q(u_usb_device_controller_s_nyet),
    .D(u_usb_device_controller_n1581),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_s_nyet_9),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/s_nyet_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/s_state_8_s2  (
    .Q(u_usb_device_controller_u_usb_packet_s_state[8]),
    .D(u_usb_device_controller_u_usb_packet_n620),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_state_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_8_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/s_state_7_s2  (
    .Q(u_usb_device_controller_u_usb_packet_s_state[7]),
    .D(u_usb_device_controller_u_usb_packet_n622),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_state_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_7_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/s_state_6_s4  (
    .Q(u_usb_device_controller_u_usb_packet_s_state[6]),
    .D(u_usb_device_controller_u_usb_packet_n624),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n615),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_6_s4 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/s_state_5_s12  (
    .Q(u_usb_device_controller_u_usb_packet_s_state[5]),
    .D(u_usb_device_controller_u_usb_packet_n626),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_state_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_5_s12 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/s_state_4_s12  (
    .Q(u_usb_device_controller_u_usb_packet_s_state[4]),
    .D(u_usb_device_controller_u_usb_packet_n628),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_state_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_4_s12 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/s_state_3_s12  (
    .Q(u_usb_device_controller_u_usb_packet_s_state[3]),
    .D(u_usb_device_controller_u_usb_packet_n630),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_state_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_3_s12 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/s_state_2_s12  (
    .Q(u_usb_device_controller_u_usb_packet_s_state[2]),
    .D(u_usb_device_controller_u_usb_packet_n632),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_state_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_2_s12 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/s_state_1_s2  (
    .Q(u_usb_device_controller_u_usb_packet_s_state[1]),
    .D(u_usb_device_controller_u_usb_packet_n633),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_n615),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_1_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_packet/s_state_0_s12  (
    .Q(u_usb_device_controller_u_usb_packet_s_state[0]),
    .D(u_usb_device_controller_u_usb_packet_n635),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_packet_s_state_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_0_s12 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_12_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[12]),
    .D(u_usb_device_controller_usb_transact_inst_n1086),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_12_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_11_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[11]),
    .D(u_usb_device_controller_usb_transact_inst_n1088),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_11_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_10_s1  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[10]),
    .D(u_usb_device_controller_usb_transact_inst_n1090),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_10_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_9_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[9]),
    .D(u_usb_device_controller_usb_transact_inst_n1091_56),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_9_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_8_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .D(u_usb_device_controller_usb_transact_inst_n1093),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_8_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_7_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[7]),
    .D(u_usb_device_controller_usb_transact_inst_n1095),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_7_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_6_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[6]),
    .D(u_usb_device_controller_usb_transact_inst_n1097),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_6_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_5_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[5]),
    .D(u_usb_device_controller_usb_transact_inst_n1099),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_5_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_4_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .D(u_usb_device_controller_usb_transact_inst_n1101),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_4_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_3_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[3]),
    .D(u_usb_device_controller_usb_transact_inst_n1103),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_3_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_2_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[2]),
    .D(u_usb_device_controller_usb_transact_inst_n1105),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_2_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_1_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[1]),
    .D(u_usb_device_controller_usb_transact_inst_n1107),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_1_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_state_0_s1  (
    .Q(u_usb_device_controller_usb_transact_inst_s_state[0]),
    .D(u_usb_device_controller_usb_transact_inst_n1109),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1091),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_state_0_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_in_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_in),
    .D(u_usb_device_controller_usb_transact_inst_n1064),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1064_23),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_in_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_out_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_out),
    .D(u_usb_device_controller_usb_transact_inst_n1066),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1064_23),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_out_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_sof_s4  (
    .Q(u_usb_device_controller_usb_transact_inst_s_sof),
    .D(u_usb_device_controller_usb_transact_inst_n1111),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_s_sof_11),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sof_s4 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_in_valid_s4  (
    .Q(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .D(u_usb_device_controller_usb_transact_inst_n1074),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1074_19),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_in_valid_s4 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_out_valid_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_out_valid),
    .D(u_usb_device_controller_usb_transact_inst_n1076),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1076_26),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_out_valid_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_sof_valid_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_sof_o_d),
    .D(u_usb_device_controller_usb_transact_inst_n1041),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_s_sof_valid),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sof_valid_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_ping_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_ping),
    .D(u_usb_device_controller_usb_transact_inst_n1070),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1064_23),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_ping_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_finished_s4  (
    .Q(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .D(u_usb_device_controller_usb_transact_inst_n1072),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1072_15),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_finished_s4 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_15_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[15]),
    .D(u_usb_device_controller_usb_transact_inst_n1118),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_wait_count_9),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_15_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_14_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[14]),
    .D(u_usb_device_controller_usb_transact_inst_n1121),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_wait_count_9),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_14_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_13_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[13]),
    .D(u_usb_device_controller_usb_transact_inst_n1124),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_wait_count_9),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_13_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_12_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[12]),
    .D(u_usb_device_controller_usb_transact_inst_n1127),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_wait_count_9),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_12_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_11_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[11]),
    .D(u_usb_device_controller_usb_transact_inst_n1130),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_wait_count_9),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_11_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_10_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[10]),
    .D(u_usb_device_controller_usb_transact_inst_n1133),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_wait_count_9),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_10_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_9_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[9]),
    .D(u_usb_device_controller_usb_transact_inst_n1136),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_wait_count_9),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_9_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_8_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[8]),
    .D(u_usb_device_controller_usb_transact_inst_n1138),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1138_41),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_8_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_7_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[7]),
    .D(u_usb_device_controller_usb_transact_inst_n1140),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1138_41),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_7_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_6_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[6]),
    .D(u_usb_device_controller_usb_transact_inst_n1142),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1138_41),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_6_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_5_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[5]),
    .D(u_usb_device_controller_usb_transact_inst_n1144),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1138_41),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_5_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_4_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[4]),
    .D(u_usb_device_controller_usb_transact_inst_n1146),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1138_41),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_4_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_3_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[3]),
    .D(u_usb_device_controller_usb_transact_inst_n1148),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1138_41),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_3_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_2_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[2]),
    .D(u_usb_device_controller_usb_transact_inst_n1150),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1138_41),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_2_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_1_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[1]),
    .D(u_usb_device_controller_usb_transact_inst_n1152),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1138_41),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_1_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/wait_count_0_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_wait_count[0]),
    .D(u_usb_device_controller_usb_transact_inst_n1154),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1138_41),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_0_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_sendpid[3]),
    .D(u_usb_device_controller_usb_transact_inst_n1157),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_s_sendpid_0),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_sendpid_2_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_sendpid[2]),
    .D(u_usb_device_controller_usb_transact_inst_n1159),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_s_sendpid_0),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_2_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_sendpid_1_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_sendpid[1]),
    .D(u_usb_device_controller_usb_transact_inst_n1161),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_n1157_23),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_1_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_transact_inst/s_sendpid_0_s2  (
    .Q(u_usb_device_controller_usb_transact_inst_s_sendpid[0]),
    .D(u_usb_device_controller_usb_transact_inst_n1163),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_transact_inst_s_sendpid_0),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_0_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_9_s2  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[9]),
    .D(u_usb_device_controller_usb_control_inst_n1672),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_9_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_8_s4  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[8]),
    .D(u_usb_device_controller_usb_control_inst_n1674),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_8_s4 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_7_s6  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[7]),
    .D(u_usb_device_controller_usb_control_inst_n1676),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_7_s6 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_6_s6  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[6]),
    .D(u_usb_device_controller_usb_control_inst_n1678),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_6_s6 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_5_s1  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[5]),
    .D(u_usb_device_controller_usb_control_inst_n1680),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_5_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_4_s6  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[4]),
    .D(u_usb_device_controller_usb_control_inst_n1682),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_4_s6 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_3_s6  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[3]),
    .D(u_usb_device_controller_usb_control_inst_n1684),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_3_s6 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_2_s6  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[2]),
    .D(u_usb_device_controller_usb_control_inst_n1686),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_2_s6 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_1_s6  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[1]),
    .D(u_usb_device_controller_usb_control_inst_n1688),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_1_s6 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_state_0_s4  (
    .Q(u_usb_device_controller_usb_control_inst_s_state[0]),
    .D(u_usb_device_controller_usb_control_inst_n1690),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_n1670),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_state_0_s4 .INIT=1'b0;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_1_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[1]),
    .D(u_usb_device_controller_usb_control_inst_n1701),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_1),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_1_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_2_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[2]),
    .D(u_usb_device_controller_usb_control_inst_n1703),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_2),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_2_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_3_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[3]),
    .D(u_usb_device_controller_usb_control_inst_n1705),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_3),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_3_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_4_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[4]),
    .D(u_usb_device_controller_usb_control_inst_n1707),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_4),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_4_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_5_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[5]),
    .D(u_usb_device_controller_usb_control_inst_n1709),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_5),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_5_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_6_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[6]),
    .D(u_usb_device_controller_usb_control_inst_n1711),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_6),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_6_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_7_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[7]),
    .D(u_usb_device_controller_usb_control_inst_n1713),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_7),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_7_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_8_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[8]),
    .D(u_usb_device_controller_usb_control_inst_n1715),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_8),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_8_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_9_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[9]),
    .D(u_usb_device_controller_usb_control_inst_n1717),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_9),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_9_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_10_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[10]),
    .D(u_usb_device_controller_usb_control_inst_n1719),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_10),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_10_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_11_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[11]),
    .D(u_usb_device_controller_usb_control_inst_n1721),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_11),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_11_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_12_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[12]),
    .D(u_usb_device_controller_usb_control_inst_n1723),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_12),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_12_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_13_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[13]),
    .D(u_usb_device_controller_usb_control_inst_n1725),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_13),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_13_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_14_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[14]),
    .D(u_usb_device_controller_usb_control_inst_n1727),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_14),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_14_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLRIN_15_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_in[15]),
    .D(u_usb_device_controller_usb_control_inst_n1729),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLRIN_15),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_15_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_1_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[1]),
    .D(u_usb_device_controller_usb_control_inst_n1731),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_1),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_1_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_2_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[2]),
    .D(u_usb_device_controller_usb_control_inst_n1733),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_2),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_2_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_3_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[3]),
    .D(u_usb_device_controller_usb_control_inst_n1735),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_3),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_3_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_4_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[4]),
    .D(u_usb_device_controller_usb_control_inst_n1737),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_4),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_4_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_5_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[5]),
    .D(u_usb_device_controller_usb_control_inst_n1739),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_5),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_5_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_6_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[6]),
    .D(u_usb_device_controller_usb_control_inst_n1741),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_6),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_6_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_7_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[7]),
    .D(u_usb_device_controller_usb_control_inst_n1743),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_7),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_7_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_8_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[8]),
    .D(u_usb_device_controller_usb_control_inst_n1745),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_8),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_8_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_9_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[9]),
    .D(u_usb_device_controller_usb_control_inst_n1747),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_9),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_9_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_10_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[10]),
    .D(u_usb_device_controller_usb_control_inst_n1749),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_10),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_10_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_11_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[11]),
    .D(u_usb_device_controller_usb_control_inst_n1751),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_11),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_11_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_12_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[12]),
    .D(u_usb_device_controller_usb_control_inst_n1753),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_12),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_12_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_13_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[13]),
    .D(u_usb_device_controller_usb_control_inst_n1755),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_13),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_13_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_14_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[14]),
    .D(u_usb_device_controller_usb_control_inst_n1757),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_14),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_14_s2 .INIT=1'b1;
  DFFSE \u_usb_device_controller/usb_control_inst/C_CLROUT_15_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_clr_out[15]),
    .D(u_usb_device_controller_usb_control_inst_n1759),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_CLROUT_15),
    .SET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_15_s2 .INIT=1'b1;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_1_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[1]),
    .D(u_usb_device_controller_usb_control_inst_n1761),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_1),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_1_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_2_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[2]),
    .D(u_usb_device_controller_usb_control_inst_n1763),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_2),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_2_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_3_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[3]),
    .D(u_usb_device_controller_usb_control_inst_n1765),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_3_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_4_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[4]),
    .D(u_usb_device_controller_usb_control_inst_n1767),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_4),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_4_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_5_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[5]),
    .D(u_usb_device_controller_usb_control_inst_n1769),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_5),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_5_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_6_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[6]),
    .D(u_usb_device_controller_usb_control_inst_n1771),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_6),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_6_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_7_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[7]),
    .D(u_usb_device_controller_usb_control_inst_n1773),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_7),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_7_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_8_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[8]),
    .D(u_usb_device_controller_usb_control_inst_n1775),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_8),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_8_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_9_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[9]),
    .D(u_usb_device_controller_usb_control_inst_n1777),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_9),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_9_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_10_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[10]),
    .D(u_usb_device_controller_usb_control_inst_n1779),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_10),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_10_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_11_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[11]),
    .D(u_usb_device_controller_usb_control_inst_n1781),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_11),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_11_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_12_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[12]),
    .D(u_usb_device_controller_usb_control_inst_n1783),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_12),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_12_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_13_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[13]),
    .D(u_usb_device_controller_usb_control_inst_n1785),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_13),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_13_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_14_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[14]),
    .D(u_usb_device_controller_usb_control_inst_n1787),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_14),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_14_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTIN_15_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[15]),
    .D(u_usb_device_controller_usb_control_inst_n1789),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTIN_15),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_15_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_1_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[1]),
    .D(u_usb_device_controller_usb_control_inst_n1791),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_1),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_1_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_2_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[2]),
    .D(u_usb_device_controller_usb_control_inst_n1793),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_2),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_2_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_3_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[3]),
    .D(u_usb_device_controller_usb_control_inst_n1795),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_3),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_3_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_4_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[4]),
    .D(u_usb_device_controller_usb_control_inst_n1797),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_4),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_4_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_5_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[5]),
    .D(u_usb_device_controller_usb_control_inst_n1799),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_5),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_5_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_6_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[6]),
    .D(u_usb_device_controller_usb_control_inst_n1801),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_6),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_6_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_7_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[7]),
    .D(u_usb_device_controller_usb_control_inst_n1803),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_7),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_7_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_8_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[8]),
    .D(u_usb_device_controller_usb_control_inst_n1805),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_8),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_8_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_9_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[9]),
    .D(u_usb_device_controller_usb_control_inst_n1807),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_9),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_9_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_10_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[10]),
    .D(u_usb_device_controller_usb_control_inst_n1809),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_10),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_10_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_11_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[11]),
    .D(u_usb_device_controller_usb_control_inst_n1811),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_11),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_11_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_12_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[12]),
    .D(u_usb_device_controller_usb_control_inst_n1813),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_12),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_12_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_13_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[13]),
    .D(u_usb_device_controller_usb_control_inst_n1815),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_13),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_13_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_14_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[14]),
    .D(u_usb_device_controller_usb_control_inst_n1817),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_14),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_14_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/C_SHLTOUT_15_s2  (
    .Q(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[15]),
    .D(u_usb_device_controller_usb_control_inst_n1819),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_C_SHLTOUT_15),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_15_s2 .INIT=1'b0;
  DFFRE \u_usb_device_controller/usb_control_inst/s_interface_set_s2  (
    .Q(u_usb_device_controller_usb_control_inst_inf_set_o_d),
    .D(u_usb_device_controller_usb_control_inst_n1629),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_usb_control_inst_s_interface_set),
    .RESET(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_interface_set_s2 .INIT=1'b0;
  ALU \u_usb_device_controller/n1473_s24  (
    .SUM(u_usb_device_controller_n1473),
    .COUT(u_usb_device_controller_n1473_28),
    .I0(VCC),
    .I1(u_usb_device_controller_s_txbuf_stop[0]),
    .I3(GND),
    .CIN(u_usb_device_controller_s_bufptr[0]) 
);
defparam \u_usb_device_controller/n1473_s24 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s25  (
    .SUM(u_usb_device_controller_n1473_29),
    .COUT(u_usb_device_controller_n1473_30),
    .I0(u_usb_device_controller_s_bufptr[1]),
    .I1(u_usb_device_controller_s_txbuf_stop[1]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_28) 
);
defparam \u_usb_device_controller/n1473_s25 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s26  (
    .SUM(u_usb_device_controller_n1473_31),
    .COUT(u_usb_device_controller_n1473_32),
    .I0(u_usb_device_controller_s_bufptr[2]),
    .I1(u_usb_device_controller_s_txbuf_stop[2]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_30) 
);
defparam \u_usb_device_controller/n1473_s26 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s27  (
    .SUM(u_usb_device_controller_n1473_33),
    .COUT(u_usb_device_controller_n1473_34),
    .I0(u_usb_device_controller_s_bufptr[3]),
    .I1(u_usb_device_controller_s_txbuf_stop[3]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_32) 
);
defparam \u_usb_device_controller/n1473_s27 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s28  (
    .SUM(u_usb_device_controller_n1473_35),
    .COUT(u_usb_device_controller_n1473_36),
    .I0(u_usb_device_controller_s_bufptr[4]),
    .I1(u_usb_device_controller_s_txbuf_stop[4]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_34) 
);
defparam \u_usb_device_controller/n1473_s28 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s29  (
    .SUM(u_usb_device_controller_n1473_37),
    .COUT(u_usb_device_controller_n1473_38),
    .I0(u_usb_device_controller_s_bufptr[5]),
    .I1(u_usb_device_controller_s_txbuf_stop[5]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_36) 
);
defparam \u_usb_device_controller/n1473_s29 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s30  (
    .SUM(u_usb_device_controller_n1473_39),
    .COUT(u_usb_device_controller_n1473_40),
    .I0(u_usb_device_controller_s_bufptr[6]),
    .I1(u_usb_device_controller_s_txbuf_stop[6]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_38) 
);
defparam \u_usb_device_controller/n1473_s30 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s31  (
    .SUM(u_usb_device_controller_n1473_41),
    .COUT(u_usb_device_controller_n1473_42),
    .I0(u_usb_device_controller_s_bufptr[7]),
    .I1(u_usb_device_controller_s_txbuf_stop[7]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_40) 
);
defparam \u_usb_device_controller/n1473_s31 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s32  (
    .SUM(u_usb_device_controller_n1473_43),
    .COUT(u_usb_device_controller_n1473_44),
    .I0(u_usb_device_controller_s_bufptr[8]),
    .I1(u_usb_device_controller_s_txbuf_stop[8]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_42) 
);
defparam \u_usb_device_controller/n1473_s32 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s33  (
    .SUM(u_usb_device_controller_n1473_45),
    .COUT(u_usb_device_controller_n1473_46),
    .I0(u_usb_device_controller_s_bufptr[9]),
    .I1(u_usb_device_controller_s_txbuf_stop[9]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_44) 
);
defparam \u_usb_device_controller/n1473_s33 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s34  (
    .SUM(u_usb_device_controller_n1473_47),
    .COUT(u_usb_device_controller_n1473_48),
    .I0(u_usb_device_controller_s_bufptr[10]),
    .I1(u_usb_device_controller_s_txbuf_stop[10]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_46) 
);
defparam \u_usb_device_controller/n1473_s34 .ALU_MODE=1;
  ALU \u_usb_device_controller/n1473_s35  (
    .SUM(u_usb_device_controller_n1473_49),
    .COUT(u_usb_device_controller_n1473_50),
    .I0(u_usb_device_controller_s_bufptr[11]),
    .I1(u_usb_device_controller_s_txbuf_stop[11]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1473_48) 
);
defparam \u_usb_device_controller/n1473_s35 .ALU_MODE=1;
  ALU \u_usb_device_controller/n2023_s  (
    .SUM(u_usb_device_controller_n2023),
    .COUT(u_usb_device_controller_n2023_2),
    .I0(u_usb_device_controller_descrom_start_0),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I3(GND),
    .CIN(GND) 
);
defparam \u_usb_device_controller/n2023_s .ALU_MODE=0;
  ALU \u_usb_device_controller/n2022_s  (
    .SUM(u_usb_device_controller_n2022),
    .COUT(u_usb_device_controller_n2022_2),
    .I0(u_usb_device_controller_descrom_start_1),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]),
    .I3(GND),
    .CIN(u_usb_device_controller_n2023_2) 
);
defparam \u_usb_device_controller/n2022_s .ALU_MODE=0;
  ALU \u_usb_device_controller/n2021_s  (
    .SUM(u_usb_device_controller_n2021),
    .COUT(u_usb_device_controller_n2021_2),
    .I0(u_usb_device_controller_descrom_start_2),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[2]),
    .I3(GND),
    .CIN(u_usb_device_controller_n2022_2) 
);
defparam \u_usb_device_controller/n2021_s .ALU_MODE=0;
  ALU \u_usb_device_controller/n2020_s  (
    .SUM(u_usb_device_controller_n2020),
    .COUT(u_usb_device_controller_n2020_2),
    .I0(u_usb_device_controller_descrom_start_3),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[3]),
    .I3(GND),
    .CIN(u_usb_device_controller_n2021_2) 
);
defparam \u_usb_device_controller/n2020_s .ALU_MODE=0;
  ALU \u_usb_device_controller/n2019_s  (
    .SUM(u_usb_device_controller_n2019),
    .COUT(u_usb_device_controller_n2019_2),
    .I0(u_usb_device_controller_descrom_start_4),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[4]),
    .I3(GND),
    .CIN(u_usb_device_controller_n2020_2) 
);
defparam \u_usb_device_controller/n2019_s .ALU_MODE=0;
  ALU \u_usb_device_controller/n2018_s  (
    .SUM(u_usb_device_controller_n2018),
    .COUT(u_usb_device_controller_n2018_2),
    .I0(u_usb_device_controller_descrom_start_5),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[5]),
    .I3(GND),
    .CIN(u_usb_device_controller_n2019_2) 
);
defparam \u_usb_device_controller/n2018_s .ALU_MODE=0;
  ALU \u_usb_device_controller/n2017_s  (
    .SUM(u_usb_device_controller_n2017),
    .COUT(u_usb_device_controller_n2017_2),
    .I0(u_usb_device_controller_descrom_start_6),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[6]),
    .I3(GND),
    .CIN(u_usb_device_controller_n2018_2) 
);
defparam \u_usb_device_controller/n2017_s .ALU_MODE=0;
  ALU \u_usb_device_controller/n2016_s  (
    .SUM(u_usb_device_controller_n2016),
    .COUT(u_usb_device_controller_n2016_2),
    .I0(u_usb_device_controller_descrom_start_7),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[7]),
    .I3(GND),
    .CIN(u_usb_device_controller_n2017_2) 
);
defparam \u_usb_device_controller/n2016_s .ALU_MODE=0;
  ALU \u_usb_device_controller/n2015_s  (
    .SUM(u_usb_device_controller_n2015),
    .COUT(u_usb_device_controller_n2015_2),
    .I0(u_usb_device_controller_descrom_start_8),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_n2016_2) 
);
defparam \u_usb_device_controller/n2015_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n240_s  (
    .SUM(u_usb_device_controller_u_usb_init_n240),
    .COUT(u_usb_device_controller_u_usb_init_n240_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[1]),
    .I1(u_usb_device_controller_u_usb_init_s_timer1[0]),
    .I3(GND),
    .CIN(GND) 
);
defparam \u_usb_device_controller/u_usb_init/n240_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n239_s  (
    .SUM(u_usb_device_controller_u_usb_init_n239),
    .COUT(u_usb_device_controller_u_usb_init_n239_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[2]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n240_2) 
);
defparam \u_usb_device_controller/u_usb_init/n239_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n238_s  (
    .SUM(u_usb_device_controller_u_usb_init_n238),
    .COUT(u_usb_device_controller_u_usb_init_n238_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[3]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n239_2) 
);
defparam \u_usb_device_controller/u_usb_init/n238_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n237_s  (
    .SUM(u_usb_device_controller_u_usb_init_n237),
    .COUT(u_usb_device_controller_u_usb_init_n237_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[4]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n238_2) 
);
defparam \u_usb_device_controller/u_usb_init/n237_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n236_s  (
    .SUM(u_usb_device_controller_u_usb_init_n236),
    .COUT(u_usb_device_controller_u_usb_init_n236_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[5]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n237_2) 
);
defparam \u_usb_device_controller/u_usb_init/n236_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n235_s  (
    .SUM(u_usb_device_controller_u_usb_init_n235),
    .COUT(u_usb_device_controller_u_usb_init_n235_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[6]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n236_2) 
);
defparam \u_usb_device_controller/u_usb_init/n235_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n234_s  (
    .SUM(u_usb_device_controller_u_usb_init_n234),
    .COUT(u_usb_device_controller_u_usb_init_n234_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[7]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n235_2) 
);
defparam \u_usb_device_controller/u_usb_init/n234_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n233_s  (
    .SUM(u_usb_device_controller_u_usb_init_n233),
    .COUT(u_usb_device_controller_u_usb_init_n233_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[8]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n234_2) 
);
defparam \u_usb_device_controller/u_usb_init/n233_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n232_s  (
    .SUM(u_usb_device_controller_u_usb_init_n232),
    .COUT(u_usb_device_controller_u_usb_init_n232_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[9]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n233_2) 
);
defparam \u_usb_device_controller/u_usb_init/n232_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n231_s  (
    .SUM(u_usb_device_controller_u_usb_init_n231),
    .COUT(u_usb_device_controller_u_usb_init_n231_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[10]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n232_2) 
);
defparam \u_usb_device_controller/u_usb_init/n231_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n230_s  (
    .SUM(u_usb_device_controller_u_usb_init_n230),
    .COUT(u_usb_device_controller_u_usb_init_n230_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[11]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n231_2) 
);
defparam \u_usb_device_controller/u_usb_init/n230_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n229_s  (
    .SUM(u_usb_device_controller_u_usb_init_n229),
    .COUT(u_usb_device_controller_u_usb_init_n229_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[12]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n230_2) 
);
defparam \u_usb_device_controller/u_usb_init/n229_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n228_s  (
    .SUM(u_usb_device_controller_u_usb_init_n228),
    .COUT(u_usb_device_controller_u_usb_init_n228_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[13]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n229_2) 
);
defparam \u_usb_device_controller/u_usb_init/n228_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n227_s  (
    .SUM(u_usb_device_controller_u_usb_init_n227),
    .COUT(u_usb_device_controller_u_usb_init_n227_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[14]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n228_2) 
);
defparam \u_usb_device_controller/u_usb_init/n227_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n226_s  (
    .SUM(u_usb_device_controller_u_usb_init_n226),
    .COUT(u_usb_device_controller_u_usb_init_n226_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[15]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n227_2) 
);
defparam \u_usb_device_controller/u_usb_init/n226_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n278_s  (
    .SUM(u_usb_device_controller_u_usb_init_n278),
    .COUT(u_usb_device_controller_u_usb_init_n278_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[1]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[0]),
    .I3(GND),
    .CIN(GND) 
);
defparam \u_usb_device_controller/u_usb_init/n278_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n277_s  (
    .SUM(u_usb_device_controller_u_usb_init_n277),
    .COUT(u_usb_device_controller_u_usb_init_n277_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[2]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n278_2) 
);
defparam \u_usb_device_controller/u_usb_init/n277_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n276_s  (
    .SUM(u_usb_device_controller_u_usb_init_n276),
    .COUT(u_usb_device_controller_u_usb_init_n276_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[3]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n277_2) 
);
defparam \u_usb_device_controller/u_usb_init/n276_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n275_s  (
    .SUM(u_usb_device_controller_u_usb_init_n275),
    .COUT(u_usb_device_controller_u_usb_init_n275_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[4]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n276_2) 
);
defparam \u_usb_device_controller/u_usb_init/n275_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n274_s  (
    .SUM(u_usb_device_controller_u_usb_init_n274),
    .COUT(u_usb_device_controller_u_usb_init_n274_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[5]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n275_2) 
);
defparam \u_usb_device_controller/u_usb_init/n274_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n273_s  (
    .SUM(u_usb_device_controller_u_usb_init_n273),
    .COUT(u_usb_device_controller_u_usb_init_n273_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[6]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n274_2) 
);
defparam \u_usb_device_controller/u_usb_init/n273_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n272_s  (
    .SUM(u_usb_device_controller_u_usb_init_n272),
    .COUT(u_usb_device_controller_u_usb_init_n272_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[7]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n273_2) 
);
defparam \u_usb_device_controller/u_usb_init/n272_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n271_s  (
    .SUM(u_usb_device_controller_u_usb_init_n271),
    .COUT(u_usb_device_controller_u_usb_init_n271_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[8]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n272_2) 
);
defparam \u_usb_device_controller/u_usb_init/n271_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n270_s  (
    .SUM(u_usb_device_controller_u_usb_init_n270),
    .COUT(u_usb_device_controller_u_usb_init_n270_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[9]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n271_2) 
);
defparam \u_usb_device_controller/u_usb_init/n270_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n269_s  (
    .SUM(u_usb_device_controller_u_usb_init_n269),
    .COUT(u_usb_device_controller_u_usb_init_n269_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[10]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n270_2) 
);
defparam \u_usb_device_controller/u_usb_init/n269_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n268_s  (
    .SUM(u_usb_device_controller_u_usb_init_n268),
    .COUT(u_usb_device_controller_u_usb_init_n268_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[11]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n269_2) 
);
defparam \u_usb_device_controller/u_usb_init/n268_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n267_s  (
    .SUM(u_usb_device_controller_u_usb_init_n267),
    .COUT(u_usb_device_controller_u_usb_init_n267_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[12]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n268_2) 
);
defparam \u_usb_device_controller/u_usb_init/n267_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n266_s  (
    .SUM(u_usb_device_controller_u_usb_init_n266),
    .COUT(u_usb_device_controller_u_usb_init_n266_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[13]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n267_2) 
);
defparam \u_usb_device_controller/u_usb_init/n266_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n265_s  (
    .SUM(u_usb_device_controller_u_usb_init_n265),
    .COUT(u_usb_device_controller_u_usb_init_n265_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[14]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n266_2) 
);
defparam \u_usb_device_controller/u_usb_init/n265_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n264_s  (
    .SUM(u_usb_device_controller_u_usb_init_n264),
    .COUT(u_usb_device_controller_u_usb_init_n264_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[15]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n265_2) 
);
defparam \u_usb_device_controller/u_usb_init/n264_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n263_s  (
    .SUM(u_usb_device_controller_u_usb_init_n263),
    .COUT(u_usb_device_controller_u_usb_init_n263_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[16]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n264_2) 
);
defparam \u_usb_device_controller/u_usb_init/n263_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n262_s  (
    .SUM(u_usb_device_controller_u_usb_init_n262),
    .COUT(u_usb_device_controller_u_usb_init_n262_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[17]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n263_2) 
);
defparam \u_usb_device_controller/u_usb_init/n262_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n261_s  (
    .SUM(u_usb_device_controller_u_usb_init_n261),
    .COUT(u_usb_device_controller_u_usb_init_n261_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[18]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n262_2) 
);
defparam \u_usb_device_controller/u_usb_init/n261_s .ALU_MODE=0;
  ALU \u_usb_device_controller/u_usb_init/n260_s  (
    .SUM(u_usb_device_controller_u_usb_init_n260),
    .COUT(u_usb_device_controller_u_usb_init_n260_2),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[19]),
    .I1(GND),
    .I3(GND),
    .CIN(u_usb_device_controller_u_usb_init_n261_2) 
);
defparam \u_usb_device_controller/u_usb_init/n260_s .ALU_MODE=0;
  DFFRE \u_usb_device_controller/isync_1_s1  (
    .Q(u_usb_device_controller_isync[1]),
    .D(u_usb_device_controller_n384),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_1),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_1_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_1_s1  (
    .Q(u_usb_device_controller_osync[1]),
    .D(u_usb_device_controller_n385),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n385_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_1_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_2_s1  (
    .Q(u_usb_device_controller_isync[2]),
    .D(u_usb_device_controller_n442),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_2),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_2_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_2_s1  (
    .Q(u_usb_device_controller_osync[2]),
    .D(u_usb_device_controller_n443),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n443_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_2_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_3_s1  (
    .Q(u_usb_device_controller_isync[3]),
    .D(u_usb_device_controller_n502),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_3),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_3_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_3_s1  (
    .Q(u_usb_device_controller_osync[3]),
    .D(u_usb_device_controller_n503),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n503_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_3_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_4_s1  (
    .Q(u_usb_device_controller_isync[4]),
    .D(u_usb_device_controller_n560),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_4),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_4_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_4_s1  (
    .Q(u_usb_device_controller_osync[4]),
    .D(u_usb_device_controller_n561),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n561_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_4_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_5_s1  (
    .Q(u_usb_device_controller_isync[5]),
    .D(u_usb_device_controller_n620),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_5),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_5_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_5_s1  (
    .Q(u_usb_device_controller_osync[5]),
    .D(u_usb_device_controller_n621),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n621_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_5_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_6_s1  (
    .Q(u_usb_device_controller_isync[6]),
    .D(u_usb_device_controller_n680),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_6_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_6_s1  (
    .Q(u_usb_device_controller_osync[6]),
    .D(u_usb_device_controller_n681),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n681_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_6_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_7_s1  (
    .Q(u_usb_device_controller_isync[7]),
    .D(u_usb_device_controller_n742),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_7),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_7_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_7_s1  (
    .Q(u_usb_device_controller_osync[7]),
    .D(u_usb_device_controller_n743),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n743_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_7_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_8_s1  (
    .Q(u_usb_device_controller_isync[8]),
    .D(u_usb_device_controller_n800),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_8),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_8_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_8_s1  (
    .Q(u_usb_device_controller_osync[8]),
    .D(u_usb_device_controller_n801),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n801_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_8_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_9_s1  (
    .Q(u_usb_device_controller_isync[9]),
    .D(u_usb_device_controller_n860),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_9),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_9_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_9_s1  (
    .Q(u_usb_device_controller_osync[9]),
    .D(u_usb_device_controller_n861),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n861_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_9_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_10_s1  (
    .Q(u_usb_device_controller_isync[10]),
    .D(u_usb_device_controller_n920),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_10),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_10_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_10_s1  (
    .Q(u_usb_device_controller_osync[10]),
    .D(u_usb_device_controller_n921),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n921_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_10_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_11_s1  (
    .Q(u_usb_device_controller_isync[11]),
    .D(u_usb_device_controller_n982),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_11),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_11_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_11_s1  (
    .Q(u_usb_device_controller_osync[11]),
    .D(u_usb_device_controller_n983),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n983_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_11_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_12_s1  (
    .Q(u_usb_device_controller_isync[12]),
    .D(u_usb_device_controller_n1042),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_12),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_12_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_12_s1  (
    .Q(u_usb_device_controller_osync[12]),
    .D(u_usb_device_controller_n1043),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n1043_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_12_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_13_s1  (
    .Q(u_usb_device_controller_isync[13]),
    .D(u_usb_device_controller_n1104),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_13),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_13_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_13_s1  (
    .Q(u_usb_device_controller_osync[13]),
    .D(u_usb_device_controller_n1105),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n1105_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_13_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_14_s1  (
    .Q(u_usb_device_controller_isync[14]),
    .D(u_usb_device_controller_n1166),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_14),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_14_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_14_s1  (
    .Q(u_usb_device_controller_osync[14]),
    .D(u_usb_device_controller_n1167),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n1167_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_14_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/isync_15_s1  (
    .Q(u_usb_device_controller_isync[15]),
    .D(u_usb_device_controller_n1230),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_isync_15),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/isync_15_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/osync_15_s1  (
    .Q(u_usb_device_controller_osync[15]),
    .D(u_usb_device_controller_n1231),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_n1231_6),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/osync_15_s1 .INIT=1'b0;
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_11_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[11]),
    .D(u_usb_device_controller_test_packet_inst_n127),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_10_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[10]),
    .D(u_usb_device_controller_test_packet_inst_n128),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_9_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[9]),
    .D(u_usb_device_controller_test_packet_inst_n129),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_8_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[8]),
    .D(u_usb_device_controller_test_packet_inst_n130),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_7_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[7]),
    .D(u_usb_device_controller_test_packet_inst_n131),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_6_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[6]),
    .D(u_usb_device_controller_test_packet_inst_n132),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_5_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[5]),
    .D(u_usb_device_controller_test_packet_inst_n133),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_4_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[4]),
    .D(u_usb_device_controller_test_packet_inst_n134),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_3_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[3]),
    .D(u_usb_device_controller_test_packet_inst_n135),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_2_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[2]),
    .D(u_usb_device_controller_test_packet_inst_n136),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_1_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[1]),
    .D(u_usb_device_controller_test_packet_inst_n137),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/cnt_0_s1  (
    .Q(u_usb_device_controller_test_packet_inst_cnt[0]),
    .D(u_usb_device_controller_test_packet_inst_n138),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_cnt_11),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_data_7_s1  (
    .Q(u_usb_device_controller_test_packet_inst_test_data_Z[7]),
    .D(u_usb_device_controller_test_packet_inst_n311),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_test_data_7),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_data_6_s1  (
    .Q(u_usb_device_controller_test_packet_inst_test_data_Z[6]),
    .D(u_usb_device_controller_test_packet_inst_n312),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_test_data_7),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_data_5_s1  (
    .Q(u_usb_device_controller_test_packet_inst_test_data_Z[5]),
    .D(u_usb_device_controller_test_packet_inst_n313),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_test_data_7),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_data_4_s1  (
    .Q(u_usb_device_controller_test_packet_inst_test_data_Z[4]),
    .D(u_usb_device_controller_test_packet_inst_n314),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_test_data_7),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_data_3_s1  (
    .Q(u_usb_device_controller_test_packet_inst_test_data_Z[3]),
    .D(u_usb_device_controller_test_packet_inst_n315),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_test_data_7),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_data_2_s1  (
    .Q(u_usb_device_controller_test_packet_inst_test_data_Z[2]),
    .D(u_usb_device_controller_test_packet_inst_n316),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_test_data_7),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_data_1_s1  (
    .Q(u_usb_device_controller_test_packet_inst_test_data_Z[1]),
    .D(u_usb_device_controller_test_packet_inst_n317),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_test_data_7),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_data_0_s1  (
    .Q(u_usb_device_controller_test_packet_inst_test_data_Z[0]),
    .D(u_usb_device_controller_test_packet_inst_n318),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_test_data_7),
    .CLEAR(reset_i_d) 
);
  DFFCE \u_usb_device_controller/test_packet_inst/test_data_val_s1  (
    .Q(u_usb_device_controller_test_packet_inst_test_dval),
    .D(u_usb_device_controller_test_packet_inst_n319),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_test_packet_inst_test_data_val),
    .CLEAR(reset_i_d) 
);
  DFFRE \u_usb_device_controller/u_usb_init/s_state_2_s1  (
    .Q(u_usb_device_controller_u_usb_init_s_state[2]),
    .D(u_usb_device_controller_u_usb_init_n215),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_state_2),
    .RESET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_2_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_state_1_s1  (
    .Q(u_usb_device_controller_u_usb_init_s_state[1]),
    .D(u_usb_device_controller_u_usb_init_n216),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_state_1),
    .RESET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_1_s1 .INIT=1'b0;
  DFFRE \u_usb_device_controller/u_usb_init/s_state_0_s1  (
    .Q(u_usb_device_controller_u_usb_init_s_state_0_4),
    .D(u_usb_device_controller_u_usb_init_n217),
    .CLK(clk_i_d),
    .CE(u_usb_device_controller_u_usb_init_s_state_0),
    .RESET(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_0_s1 .INIT=1'b0;
  ALU \u_usb_device_controller/n1454_s0  (
    .SUM(u_usb_device_controller_n1454),
    .COUT(u_usb_device_controller_n1454_3),
    .I0(u_usb_device_controller_s_bufptr[0]),
    .I1(u_usb_device_controller_s_txbuf_stop[0]),
    .I3(GND),
    .CIN(GND) 
);
defparam \u_usb_device_controller/n1454_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1455_s0  (
    .SUM(u_usb_device_controller_n1455),
    .COUT(u_usb_device_controller_n1455_3),
    .I0(u_usb_device_controller_s_bufptr[1]),
    .I1(u_usb_device_controller_s_txbuf_stop[1]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1454_3) 
);
defparam \u_usb_device_controller/n1455_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1456_s0  (
    .SUM(u_usb_device_controller_n1456),
    .COUT(u_usb_device_controller_n1456_3),
    .I0(u_usb_device_controller_s_bufptr[2]),
    .I1(u_usb_device_controller_s_txbuf_stop[2]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1455_3) 
);
defparam \u_usb_device_controller/n1456_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1457_s0  (
    .SUM(u_usb_device_controller_n1457),
    .COUT(u_usb_device_controller_n1457_3),
    .I0(u_usb_device_controller_s_bufptr[3]),
    .I1(u_usb_device_controller_s_txbuf_stop[3]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1456_3) 
);
defparam \u_usb_device_controller/n1457_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1458_s0  (
    .SUM(u_usb_device_controller_n1458),
    .COUT(u_usb_device_controller_n1458_3),
    .I0(u_usb_device_controller_s_bufptr[4]),
    .I1(u_usb_device_controller_s_txbuf_stop[4]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1457_3) 
);
defparam \u_usb_device_controller/n1458_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1459_s0  (
    .SUM(u_usb_device_controller_n1459),
    .COUT(u_usb_device_controller_n1459_3),
    .I0(u_usb_device_controller_s_bufptr[5]),
    .I1(u_usb_device_controller_s_txbuf_stop[5]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1458_3) 
);
defparam \u_usb_device_controller/n1459_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1460_s0  (
    .SUM(u_usb_device_controller_n1460),
    .COUT(u_usb_device_controller_n1460_3),
    .I0(u_usb_device_controller_s_bufptr[6]),
    .I1(u_usb_device_controller_s_txbuf_stop[6]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1459_3) 
);
defparam \u_usb_device_controller/n1460_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1461_s0  (
    .SUM(u_usb_device_controller_n1461),
    .COUT(u_usb_device_controller_n1461_3),
    .I0(u_usb_device_controller_s_bufptr[7]),
    .I1(u_usb_device_controller_s_txbuf_stop[7]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1460_3) 
);
defparam \u_usb_device_controller/n1461_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1462_s0  (
    .SUM(u_usb_device_controller_n1462),
    .COUT(u_usb_device_controller_n1462_3),
    .I0(u_usb_device_controller_s_bufptr[8]),
    .I1(u_usb_device_controller_s_txbuf_stop[8]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1461_3) 
);
defparam \u_usb_device_controller/n1462_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1463_s0  (
    .SUM(u_usb_device_controller_n1463),
    .COUT(u_usb_device_controller_n1463_3),
    .I0(u_usb_device_controller_s_bufptr[9]),
    .I1(u_usb_device_controller_s_txbuf_stop[9]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1462_3) 
);
defparam \u_usb_device_controller/n1463_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1464_s0  (
    .SUM(u_usb_device_controller_n1464),
    .COUT(u_usb_device_controller_n1464_3),
    .I0(u_usb_device_controller_s_bufptr[10]),
    .I1(u_usb_device_controller_s_txbuf_stop[10]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1463_3) 
);
defparam \u_usb_device_controller/n1464_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/n1465_s0  (
    .SUM(u_usb_device_controller_n1465),
    .COUT(u_usb_device_controller_n1465_3),
    .I0(u_usb_device_controller_s_bufptr[11]),
    .I1(u_usb_device_controller_s_txbuf_stop[11]),
    .I3(GND),
    .CIN(u_usb_device_controller_n1464_3) 
);
defparam \u_usb_device_controller/n1465_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_transact_inst/n156_s0  (
    .SUM(u_usb_device_controller_usb_transact_inst_n156),
    .COUT(u_usb_device_controller_usb_transact_inst_n156_3),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_addr[0]),
    .I3(GND),
    .CIN(GND) 
);
defparam \u_usb_device_controller/usb_transact_inst/n156_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_transact_inst/n157_s0  (
    .SUM(u_usb_device_controller_usb_transact_inst_n157),
    .COUT(u_usb_device_controller_usb_transact_inst_n157_3),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_addr[1]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_transact_inst_n156_3) 
);
defparam \u_usb_device_controller/usb_transact_inst/n157_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_transact_inst/n158_s0  (
    .SUM(u_usb_device_controller_usb_transact_inst_n158),
    .COUT(u_usb_device_controller_usb_transact_inst_n158_3),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_addr[2]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_transact_inst_n157_3) 
);
defparam \u_usb_device_controller/usb_transact_inst/n158_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_transact_inst/n159_s0  (
    .SUM(u_usb_device_controller_usb_transact_inst_n159),
    .COUT(u_usb_device_controller_usb_transact_inst_n159_3),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_addr[3]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_transact_inst_n158_3) 
);
defparam \u_usb_device_controller/usb_transact_inst/n159_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_transact_inst/n160_s0  (
    .SUM(u_usb_device_controller_usb_transact_inst_n160),
    .COUT(u_usb_device_controller_usb_transact_inst_n160_3),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_addr[4]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_transact_inst_n159_3) 
);
defparam \u_usb_device_controller/usb_transact_inst/n160_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_transact_inst/n161_s0  (
    .SUM(u_usb_device_controller_usb_transact_inst_n161),
    .COUT(u_usb_device_controller_usb_transact_inst_n161_3),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_addr[5]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_transact_inst_n160_3) 
);
defparam \u_usb_device_controller/usb_transact_inst/n161_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_transact_inst/n162_s0  (
    .SUM(u_usb_device_controller_usb_transact_inst_n162),
    .COUT(u_usb_device_controller_usb_transact_inst_n162_3),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_addr[6]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_transact_inst_n161_3) 
);
defparam \u_usb_device_controller/usb_transact_inst/n162_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1467_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1467),
    .COUT(u_usb_device_controller_usb_control_inst_n1467_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I1(u_usb_device_controller_usbc_dsclen_0),
    .I3(GND),
    .CIN(GND) 
);
defparam \u_usb_device_controller/usb_control_inst/n1467_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1468_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1468),
    .COUT(u_usb_device_controller_usb_control_inst_n1468_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]),
    .I1(u_usb_device_controller_usbc_dsclen_1),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1467_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1468_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1469_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1469),
    .COUT(u_usb_device_controller_usb_control_inst_n1469_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[2]),
    .I1(u_usb_device_controller_usbc_dsclen_2),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1468_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1469_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1470_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1470),
    .COUT(u_usb_device_controller_usb_control_inst_n1470_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[3]),
    .I1(u_usb_device_controller_usbc_dsclen_3),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1469_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1470_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1471_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1471),
    .COUT(u_usb_device_controller_usb_control_inst_n1471_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[4]),
    .I1(u_usb_device_controller_usbc_dsclen_4),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1470_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1471_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1472_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1472),
    .COUT(u_usb_device_controller_usb_control_inst_n1472_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[5]),
    .I1(u_usb_device_controller_usbc_dsclen_5),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1471_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1472_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1473_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1473),
    .COUT(u_usb_device_controller_usb_control_inst_n1473_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[6]),
    .I1(u_usb_device_controller_usbc_dsclen_6),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1472_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1473_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1474_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1474),
    .COUT(u_usb_device_controller_usb_control_inst_n1474_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[7]),
    .I1(u_usb_device_controller_usbc_dsclen_7),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1473_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1474_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1476_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1476),
    .COUT(u_usb_device_controller_usb_control_inst_n1476_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen[0]),
    .I3(GND),
    .CIN(GND) 
);
defparam \u_usb_device_controller/usb_control_inst/n1476_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1477_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1477),
    .COUT(u_usb_device_controller_usb_control_inst_n1477_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen[1]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1476_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1477_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1478_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1478),
    .COUT(u_usb_device_controller_usb_control_inst_n1478_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[2]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen[2]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1477_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1478_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1479_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1479),
    .COUT(u_usb_device_controller_usb_control_inst_n1479_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[3]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen[3]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1478_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1479_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1480_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1480),
    .COUT(u_usb_device_controller_usb_control_inst_n1480_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[4]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen[4]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1479_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1480_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1481_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1481),
    .COUT(u_usb_device_controller_usb_control_inst_n1481_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[5]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen[5]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1480_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1481_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1482_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1482),
    .COUT(u_usb_device_controller_usb_control_inst_n1482_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen[6]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1481_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1482_s0 .ALU_MODE=3;
  ALU \u_usb_device_controller/usb_control_inst/n1483_s0  (
    .SUM(u_usb_device_controller_usb_control_inst_n1483),
    .COUT(u_usb_device_controller_usb_control_inst_n1483_3),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[7]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen[7]),
    .I3(GND),
    .CIN(u_usb_device_controller_usb_control_inst_n1482_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1483_s0 .ALU_MODE=3;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s43  (
    .F(u_usb_device_controller_usb_control_inst_n611),
    .I0(u_usb_device_controller_halt_out[2]),
    .I1(u_usb_device_controller_halt_in[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s43 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s44  (
    .F(u_usb_device_controller_usb_control_inst_n613),
    .I0(u_usb_device_controller_halt_out[3]),
    .I1(u_usb_device_controller_halt_in[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s44 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s45  (
    .F(u_usb_device_controller_usb_control_inst_n615),
    .I0(u_usb_device_controller_halt_out[4]),
    .I1(u_usb_device_controller_halt_in[4]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s45 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s46  (
    .F(u_usb_device_controller_usb_control_inst_n617),
    .I0(u_usb_device_controller_halt_out[5]),
    .I1(u_usb_device_controller_halt_in[5]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s46 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s47  (
    .F(u_usb_device_controller_usb_control_inst_n619),
    .I0(u_usb_device_controller_halt_out[6]),
    .I1(u_usb_device_controller_halt_in[6]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s47 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s48  (
    .F(u_usb_device_controller_usb_control_inst_n621),
    .I0(u_usb_device_controller_halt_out[7]),
    .I1(u_usb_device_controller_halt_in[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s48 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s49  (
    .F(u_usb_device_controller_usb_control_inst_n623),
    .I0(u_usb_device_controller_halt_out[8]),
    .I1(u_usb_device_controller_halt_in[8]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s49 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s50  (
    .F(u_usb_device_controller_usb_control_inst_n625),
    .I0(u_usb_device_controller_halt_out[9]),
    .I1(u_usb_device_controller_halt_in[9]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s50 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s51  (
    .F(u_usb_device_controller_usb_control_inst_n627),
    .I0(u_usb_device_controller_halt_out[10]),
    .I1(u_usb_device_controller_halt_in[10]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s51 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s52  (
    .F(u_usb_device_controller_usb_control_inst_n629),
    .I0(u_usb_device_controller_halt_out[11]),
    .I1(u_usb_device_controller_halt_in[11]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s52 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s53  (
    .F(u_usb_device_controller_usb_control_inst_n631),
    .I0(u_usb_device_controller_halt_out[12]),
    .I1(u_usb_device_controller_halt_in[12]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s53 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s54  (
    .F(u_usb_device_controller_usb_control_inst_n633),
    .I0(u_usb_device_controller_halt_out[13]),
    .I1(u_usb_device_controller_halt_in[13]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s54 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s55  (
    .F(u_usb_device_controller_usb_control_inst_n635),
    .I0(u_usb_device_controller_halt_out[14]),
    .I1(u_usb_device_controller_halt_in[14]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s55 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n645_s56  (
    .F(u_usb_device_controller_usb_control_inst_n637),
    .I0(u_usb_device_controller_halt_out[15]),
    .I1(u_usb_device_controller_halt_in[15]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n645_s56 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1241_s54  (
    .F(u_usb_device_controller_n1241_39),
    .I0(u_usb_device_controller_halt_out[4]),
    .I1(u_usb_device_controller_halt_out[5]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1241_s54 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1241_s55  (
    .F(u_usb_device_controller_n1241_40),
    .I0(u_usb_device_controller_halt_out[6]),
    .I1(u_usb_device_controller_halt_out[7]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1241_s55 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1241_s56  (
    .F(u_usb_device_controller_n1241_41),
    .I0(u_usb_device_controller_halt_out[8]),
    .I1(u_usb_device_controller_halt_out[9]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1241_s56 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1241_s57  (
    .F(u_usb_device_controller_n1241_42),
    .I0(u_usb_device_controller_halt_out[10]),
    .I1(u_usb_device_controller_halt_out[11]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1241_s57 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1241_s58  (
    .F(u_usb_device_controller_n1241_43),
    .I0(u_usb_device_controller_halt_out[12]),
    .I1(u_usb_device_controller_halt_out[13]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1241_s58 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1241_s59  (
    .F(u_usb_device_controller_n1241_44),
    .I0(u_usb_device_controller_halt_out[14]),
    .I1(u_usb_device_controller_halt_out[15]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1241_s59 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1242_s54  (
    .F(u_usb_device_controller_n1242_39),
    .I0(u_usb_device_controller_halt_in[4]),
    .I1(u_usb_device_controller_halt_in[5]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1242_s54 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1242_s55  (
    .F(u_usb_device_controller_n1242_40),
    .I0(u_usb_device_controller_halt_in[6]),
    .I1(u_usb_device_controller_halt_in[7]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1242_s55 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1242_s56  (
    .F(u_usb_device_controller_n1242_41),
    .I0(u_usb_device_controller_halt_in[8]),
    .I1(u_usb_device_controller_halt_in[9]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1242_s56 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1242_s57  (
    .F(u_usb_device_controller_n1242_42),
    .I0(u_usb_device_controller_halt_in[10]),
    .I1(u_usb_device_controller_halt_in[11]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1242_s57 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1242_s58  (
    .F(u_usb_device_controller_n1242_43),
    .I0(u_usb_device_controller_halt_in[12]),
    .I1(u_usb_device_controller_halt_in[13]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1242_s58 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1242_s59  (
    .F(u_usb_device_controller_n1242_44),
    .I0(u_usb_device_controller_halt_in[14]),
    .I1(u_usb_device_controller_halt_in[15]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1242_s59 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1243_s54  (
    .F(u_usb_device_controller_n1243_39),
    .I0(u_usb_device_controller_osync[4]),
    .I1(u_usb_device_controller_osync[5]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1243_s54 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1243_s55  (
    .F(u_usb_device_controller_n1243_40),
    .I0(u_usb_device_controller_osync[6]),
    .I1(u_usb_device_controller_osync[7]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1243_s55 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1243_s56  (
    .F(u_usb_device_controller_n1243_41),
    .I0(u_usb_device_controller_osync[8]),
    .I1(u_usb_device_controller_osync[9]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1243_s56 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1243_s57  (
    .F(u_usb_device_controller_n1243_42),
    .I0(u_usb_device_controller_osync[10]),
    .I1(u_usb_device_controller_osync[11]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1243_s57 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1243_s58  (
    .F(u_usb_device_controller_n1243_43),
    .I0(u_usb_device_controller_osync[12]),
    .I1(u_usb_device_controller_osync[13]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1243_s58 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1243_s59  (
    .F(u_usb_device_controller_n1243_44),
    .I0(u_usb_device_controller_osync[14]),
    .I1(u_usb_device_controller_osync[15]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1243_s59 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1244_s54  (
    .F(u_usb_device_controller_n1244_39),
    .I0(u_usb_device_controller_isync[4]),
    .I1(u_usb_device_controller_isync[5]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1244_s54 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1244_s55  (
    .F(u_usb_device_controller_n1244_40),
    .I0(u_usb_device_controller_isync[6]),
    .I1(u_usb_device_controller_isync[7]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1244_s55 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1244_s56  (
    .F(u_usb_device_controller_n1244_41),
    .I0(u_usb_device_controller_isync[8]),
    .I1(u_usb_device_controller_isync[9]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1244_s56 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1244_s57  (
    .F(u_usb_device_controller_n1244_42),
    .I0(u_usb_device_controller_isync[10]),
    .I1(u_usb_device_controller_isync[11]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1244_s57 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1244_s58  (
    .F(u_usb_device_controller_n1244_43),
    .I0(u_usb_device_controller_isync[12]),
    .I1(u_usb_device_controller_isync[13]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1244_s58 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1244_s59  (
    .F(u_usb_device_controller_n1244_44),
    .I0(u_usb_device_controller_isync[14]),
    .I1(u_usb_device_controller_isync[15]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1244_s59 .INIT=8'hCA;
  MUX2_LUT5 \u_usb_device_controller/usb_control_inst/n645_s24  (
    .O(u_usb_device_controller_usb_control_inst_n645),
    .I0(u_usb_device_controller_usb_control_inst_n611),
    .I1(u_usb_device_controller_usb_control_inst_n613),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
  MUX2_LUT5 \u_usb_device_controller/usb_control_inst/n645_s37  (
    .O(u_usb_device_controller_usb_control_inst_n645_33),
    .I0(u_usb_device_controller_usb_control_inst_n615),
    .I1(u_usb_device_controller_usb_control_inst_n617),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
  MUX2_LUT5 \u_usb_device_controller/usb_control_inst/n645_s38  (
    .O(u_usb_device_controller_usb_control_inst_n645_35),
    .I0(u_usb_device_controller_usb_control_inst_n619),
    .I1(u_usb_device_controller_usb_control_inst_n621),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
  MUX2_LUT5 \u_usb_device_controller/usb_control_inst/n645_s39  (
    .O(u_usb_device_controller_usb_control_inst_n645_37),
    .I0(u_usb_device_controller_usb_control_inst_n623),
    .I1(u_usb_device_controller_usb_control_inst_n625),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
  MUX2_LUT5 \u_usb_device_controller/usb_control_inst/n645_s40  (
    .O(u_usb_device_controller_usb_control_inst_n645_39),
    .I0(u_usb_device_controller_usb_control_inst_n627),
    .I1(u_usb_device_controller_usb_control_inst_n629),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
  MUX2_LUT5 \u_usb_device_controller/usb_control_inst/n645_s41  (
    .O(u_usb_device_controller_usb_control_inst_n645_41),
    .I0(u_usb_device_controller_usb_control_inst_n631),
    .I1(u_usb_device_controller_usb_control_inst_n633),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
  MUX2_LUT5 \u_usb_device_controller/usb_control_inst/n645_s42  (
    .O(u_usb_device_controller_usb_control_inst_n645_43),
    .I0(u_usb_device_controller_usb_control_inst_n635),
    .I1(u_usb_device_controller_usb_control_inst_n637),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1241_s53  (
    .O(u_usb_device_controller_n1241_46),
    .I0(u_usb_device_controller_n1241_39),
    .I1(u_usb_device_controller_n1241_40),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1241_s50  (
    .O(u_usb_device_controller_n1241_48),
    .I0(u_usb_device_controller_n1241_41),
    .I1(u_usb_device_controller_n1241_42),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1241_s51  (
    .O(u_usb_device_controller_n1241_50),
    .I0(u_usb_device_controller_n1241_43),
    .I1(u_usb_device_controller_n1241_44),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1242_s53  (
    .O(u_usb_device_controller_n1242_46),
    .I0(u_usb_device_controller_n1242_39),
    .I1(u_usb_device_controller_n1242_40),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1242_s50  (
    .O(u_usb_device_controller_n1242_48),
    .I0(u_usb_device_controller_n1242_41),
    .I1(u_usb_device_controller_n1242_42),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1242_s51  (
    .O(u_usb_device_controller_n1242_50),
    .I0(u_usb_device_controller_n1242_43),
    .I1(u_usb_device_controller_n1242_44),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1243_s53  (
    .O(u_usb_device_controller_n1243_46),
    .I0(u_usb_device_controller_n1243_39),
    .I1(u_usb_device_controller_n1243_40),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1243_s50  (
    .O(u_usb_device_controller_n1243_48),
    .I0(u_usb_device_controller_n1243_41),
    .I1(u_usb_device_controller_n1243_42),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1243_s51  (
    .O(u_usb_device_controller_n1243_50),
    .I0(u_usb_device_controller_n1243_43),
    .I1(u_usb_device_controller_n1243_44),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1244_s53  (
    .O(u_usb_device_controller_n1244_46),
    .I0(u_usb_device_controller_n1244_39),
    .I1(u_usb_device_controller_n1244_40),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1244_s50  (
    .O(u_usb_device_controller_n1244_48),
    .I0(u_usb_device_controller_n1244_41),
    .I1(u_usb_device_controller_n1244_42),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1244_s51  (
    .O(u_usb_device_controller_n1244_50),
    .I0(u_usb_device_controller_n1244_43),
    .I1(u_usb_device_controller_n1244_44),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT6 \u_usb_device_controller/n1241_s49  (
    .O(u_usb_device_controller_n1241_52),
    .I0(u_usb_device_controller_n1241_48),
    .I1(u_usb_device_controller_n1241_50),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
  MUX2_LUT6 \u_usb_device_controller/n1242_s49  (
    .O(u_usb_device_controller_n1242_52),
    .I0(u_usb_device_controller_n1242_48),
    .I1(u_usb_device_controller_n1242_50),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
  MUX2_LUT6 \u_usb_device_controller/n1243_s49  (
    .O(u_usb_device_controller_n1243_52),
    .I0(u_usb_device_controller_n1243_48),
    .I1(u_usb_device_controller_n1243_50),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
  MUX2_LUT6 \u_usb_device_controller/n1244_s49  (
    .O(u_usb_device_controller_n1244_52),
    .I0(u_usb_device_controller_n1244_48),
    .I1(u_usb_device_controller_n1244_50),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
  MUX2_LUT6 \u_usb_device_controller/usb_control_inst/n645_s31  (
    .O(u_usb_device_controller_usb_control_inst_n645_45),
    .I0(u_usb_device_controller_usb_control_inst_n645_33),
    .I1(u_usb_device_controller_usb_control_inst_n645_35),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]) 
);
  MUX2_LUT6 \u_usb_device_controller/usb_control_inst/n645_s35  (
    .O(u_usb_device_controller_usb_control_inst_n645_47),
    .I0(u_usb_device_controller_usb_control_inst_n645_37),
    .I1(u_usb_device_controller_usb_control_inst_n645_39),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]) 
);
  MUX2_LUT6 \u_usb_device_controller/usb_control_inst/n645_s36  (
    .O(u_usb_device_controller_usb_control_inst_n645_49),
    .I0(u_usb_device_controller_usb_control_inst_n645_41),
    .I1(u_usb_device_controller_usb_control_inst_n645_43),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]) 
);
  MUX2_LUT7 \u_usb_device_controller/usb_control_inst/n645_s34  (
    .O(u_usb_device_controller_usb_control_inst_n645_51),
    .I0(u_usb_device_controller_usb_control_inst_n645_47),
    .I1(u_usb_device_controller_usb_control_inst_n645_49),
    .S0(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1241_s52  (
    .O(u_usb_device_controller_n1241_54),
    .I0(u_usb_device_controller_n1241_62),
    .I1(u_usb_device_controller_n1241_60),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1242_s52  (
    .O(u_usb_device_controller_n1242_54),
    .I0(u_usb_device_controller_n1242_62),
    .I1(u_usb_device_controller_n1242_60),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1243_s52  (
    .O(u_usb_device_controller_n1243_54),
    .I0(u_usb_device_controller_n1243_62),
    .I1(u_usb_device_controller_n1243_60),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT5 \u_usb_device_controller/n1244_s52  (
    .O(u_usb_device_controller_n1244_54),
    .I0(u_usb_device_controller_n1244_62),
    .I1(u_usb_device_controller_n1244_60),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]) 
);
  MUX2_LUT6 \u_usb_device_controller/n1241_s48  (
    .O(u_usb_device_controller_n1241_56),
    .I0(u_usb_device_controller_n1241_54),
    .I1(u_usb_device_controller_n1241_46),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
  MUX2_LUT6 \u_usb_device_controller/n1242_s48  (
    .O(u_usb_device_controller_n1242_56),
    .I0(u_usb_device_controller_n1242_54),
    .I1(u_usb_device_controller_n1242_46),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
  MUX2_LUT6 \u_usb_device_controller/n1243_s48  (
    .O(u_usb_device_controller_n1243_56),
    .I0(u_usb_device_controller_n1243_54),
    .I1(u_usb_device_controller_n1243_46),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
  MUX2_LUT6 \u_usb_device_controller/n1244_s48  (
    .O(u_usb_device_controller_n1244_56),
    .I0(u_usb_device_controller_n1244_54),
    .I1(u_usb_device_controller_n1244_46),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
  MUX2_LUT7 \u_usb_device_controller/n1241_s45  (
    .O(u_usb_device_controller_n1241),
    .I0(u_usb_device_controller_n1241_56),
    .I1(u_usb_device_controller_n1241_52),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
  MUX2_LUT7 \u_usb_device_controller/n1242_s45  (
    .O(u_usb_device_controller_n1242),
    .I0(u_usb_device_controller_n1242_56),
    .I1(u_usb_device_controller_n1242_52),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
  MUX2_LUT7 \u_usb_device_controller/n1243_s45  (
    .O(u_usb_device_controller_n1243),
    .I0(u_usb_device_controller_n1243_56),
    .I1(u_usb_device_controller_n1243_52),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
  MUX2_LUT7 \u_usb_device_controller/n1244_s45  (
    .O(u_usb_device_controller_n1244),
    .I0(u_usb_device_controller_n1244_56),
    .I1(u_usb_device_controller_n1244_52),
    .S0(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
  LUT3 \u_usb_device_controller/utmi_dataout_o_d_0_s  (
    .F(u_usb_device_controller_utmi_dataout_o_d[0]),
    .I0(u_usb_device_controller_utmi_dataout_o_d_0),
    .I1(u_usb_device_controller_u_usb_packet_usbp_dataout_o[0]),
    .I2(u_usb_device_controller_test_packet_inst_test_en_dly_Z) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_0_s .INIT=8'hAC;
  LUT4 \u_usb_device_controller/utmi_txvalid_o_d_s  (
    .F(u_usb_device_controller_utmi_txvalid_o_d),
    .I0(u_usb_device_controller_test_packet_inst_test_dval),
    .I1(u_usb_device_controller_u_usb_packet_usbp_txvalid_o),
    .I2(u_usb_device_controller_utmi_txvalid_o_d_6),
    .I3(u_usb_device_controller_utmi_txvalid_o_d_8) 
);
defparam \u_usb_device_controller/utmi_txvalid_o_d_s .INIT=16'hACFF;
  LUT2 \u_usb_device_controller/n2219_s0  (
    .F(u_usb_device_controller_n2219),
    .I0(reset_i_d),
    .I1(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/n2219_s0 .INIT=4'hE;
  LUT3 \u_usb_device_controller/n384_s2  (
    .F(u_usb_device_controller_n384),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[1]),
    .I1(u_usb_device_controller_isync[1]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n384_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n385_s1  (
    .F(u_usb_device_controller_n385),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[1]),
    .I1(u_usb_device_controller_osync[1]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n385_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n442_s2  (
    .F(u_usb_device_controller_n442),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[2]),
    .I1(u_usb_device_controller_isync[2]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n442_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n443_s1  (
    .F(u_usb_device_controller_n443),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[2]),
    .I1(u_usb_device_controller_osync[2]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n443_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n502_s2  (
    .F(u_usb_device_controller_n502),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[3]),
    .I1(u_usb_device_controller_isync[3]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n502_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n503_s1  (
    .F(u_usb_device_controller_n503),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[3]),
    .I1(u_usb_device_controller_osync[3]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n503_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n560_s2  (
    .F(u_usb_device_controller_n560),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[4]),
    .I1(u_usb_device_controller_isync[4]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n560_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n561_s1  (
    .F(u_usb_device_controller_n561),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[4]),
    .I1(u_usb_device_controller_osync[4]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n561_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n620_s2  (
    .F(u_usb_device_controller_n620),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[5]),
    .I1(u_usb_device_controller_isync[5]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n620_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n621_s1  (
    .F(u_usb_device_controller_n621),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[5]),
    .I1(u_usb_device_controller_osync[5]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n621_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n680_s2  (
    .F(u_usb_device_controller_n680),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[6]),
    .I1(u_usb_device_controller_isync[6]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n680_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n681_s1  (
    .F(u_usb_device_controller_n681),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[6]),
    .I1(u_usb_device_controller_osync[6]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n681_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n742_s2  (
    .F(u_usb_device_controller_n742),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[7]),
    .I1(u_usb_device_controller_isync[7]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n742_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n743_s1  (
    .F(u_usb_device_controller_n743),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[7]),
    .I1(u_usb_device_controller_osync[7]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n743_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n800_s2  (
    .F(u_usb_device_controller_n800),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[8]),
    .I1(u_usb_device_controller_isync[8]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n800_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n801_s1  (
    .F(u_usb_device_controller_n801),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[8]),
    .I1(u_usb_device_controller_osync[8]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n801_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n860_s2  (
    .F(u_usb_device_controller_n860),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[9]),
    .I1(u_usb_device_controller_isync[9]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n860_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n861_s1  (
    .F(u_usb_device_controller_n861),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[9]),
    .I1(u_usb_device_controller_osync[9]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n861_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n920_s2  (
    .F(u_usb_device_controller_n920),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[10]),
    .I1(u_usb_device_controller_isync[10]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n920_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n921_s1  (
    .F(u_usb_device_controller_n921),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[10]),
    .I1(u_usb_device_controller_osync[10]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n921_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n982_s2  (
    .F(u_usb_device_controller_n982),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[11]),
    .I1(u_usb_device_controller_isync[11]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n982_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n983_s1  (
    .F(u_usb_device_controller_n983),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[11]),
    .I1(u_usb_device_controller_osync[11]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n983_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n1042_s2  (
    .F(u_usb_device_controller_n1042),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[12]),
    .I1(u_usb_device_controller_isync[12]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1042_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n1043_s1  (
    .F(u_usb_device_controller_n1043),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[12]),
    .I1(u_usb_device_controller_osync[12]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1043_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n1104_s2  (
    .F(u_usb_device_controller_n1104),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[13]),
    .I1(u_usb_device_controller_isync[13]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1104_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n1105_s1  (
    .F(u_usb_device_controller_n1105),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[13]),
    .I1(u_usb_device_controller_osync[13]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1105_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n1166_s2  (
    .F(u_usb_device_controller_n1166),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[14]),
    .I1(u_usb_device_controller_isync[14]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1166_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n1167_s1  (
    .F(u_usb_device_controller_n1167),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[14]),
    .I1(u_usb_device_controller_osync[14]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1167_s1 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n1230_s2  (
    .F(u_usb_device_controller_n1230),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_in[15]),
    .I1(u_usb_device_controller_isync[15]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1230_s2 .INIT=8'h43;
  LUT3 \u_usb_device_controller/n1231_s1  (
    .F(u_usb_device_controller_n1231),
    .I0(u_usb_device_controller_usb_control_inst_usbc_clr_out[15]),
    .I1(u_usb_device_controller_osync[15]),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1231_s1 .INIT=8'h43;
  LUT4 \u_usb_device_controller/n2339_s0  (
    .F(u_usb_device_controller_n2339),
    .I0(u_usb_device_controller_n2339_4),
    .I1(txdat_len_i_d[10]),
    .I2(txdat_len_i_d[11]),
    .I3(reset_i_d) 
);
defparam \u_usb_device_controller/n2339_s0 .INIT=16'hFFF4;
  LUT4 \u_usb_device_controller/txpktfin_o_d_s  (
    .F(u_usb_device_controller_txpktfin_o_d),
    .I0(u_usb_device_controller_cur_state[1]),
    .I1(u_usb_device_controller_cur_state[0]),
    .I2(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I3(u_usb_device_controller_rxact_o_d_3) 
);
defparam \u_usb_device_controller/txpktfin_o_d_s .INIT=16'h4000;
  LUT3 \u_usb_device_controller/n2025_s0  (
    .F(u_usb_device_controller_n2025),
    .I0(desc_oscfg_addr_i_d[8]),
    .I1(u_usb_device_controller_n2015),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2025_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/n2026_s0  (
    .F(u_usb_device_controller_n2026),
    .I0(desc_oscfg_addr_i_d[7]),
    .I1(u_usb_device_controller_n2016),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2026_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/n2027_s0  (
    .F(u_usb_device_controller_n2027),
    .I0(desc_oscfg_addr_i_d[6]),
    .I1(u_usb_device_controller_n2017),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2027_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/n2028_s0  (
    .F(u_usb_device_controller_n2028),
    .I0(desc_oscfg_addr_i_d[5]),
    .I1(u_usb_device_controller_n2018),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2028_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/n2029_s0  (
    .F(u_usb_device_controller_n2029),
    .I0(desc_oscfg_addr_i_d[4]),
    .I1(u_usb_device_controller_n2019),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2029_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/n2030_s0  (
    .F(u_usb_device_controller_n2030),
    .I0(desc_oscfg_addr_i_d[3]),
    .I1(u_usb_device_controller_n2020),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2030_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/n2031_s0  (
    .F(u_usb_device_controller_n2031),
    .I0(desc_oscfg_addr_i_d[2]),
    .I1(u_usb_device_controller_n2021),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2031_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/n2032_s0  (
    .F(u_usb_device_controller_n2032),
    .I0(desc_oscfg_addr_i_d[1]),
    .I1(u_usb_device_controller_n2022),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2032_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/n2033_s0  (
    .F(u_usb_device_controller_n2033),
    .I0(desc_oscfg_addr_i_d[0]),
    .I1(u_usb_device_controller_n2023),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2033_s0 .INIT=8'hAC;
  LUT4 \u_usb_device_controller/test_packet_inst/n127_s2  (
    .F(u_usb_device_controller_test_packet_inst_n127),
    .I0(u_usb_device_controller_test_packet_inst_cnt[10]),
    .I1(u_usb_device_controller_test_packet_inst_n127_6),
    .I2(u_usb_device_controller_test_packet_inst_cnt[11]),
    .I3(u_usb_device_controller_test_packet_inst_n127_7) 
);
defparam \u_usb_device_controller/test_packet_inst/n127_s2 .INIT=16'hF800;
  LUT3 \u_usb_device_controller/test_packet_inst/n128_s2  (
    .F(u_usb_device_controller_test_packet_inst_n128),
    .I0(u_usb_device_controller_test_packet_inst_cnt[10]),
    .I1(u_usb_device_controller_test_packet_inst_n127_6),
    .I2(u_usb_device_controller_test_packet_inst_n127_7) 
);
defparam \u_usb_device_controller/test_packet_inst/n128_s2 .INIT=8'h60;
  LUT4 \u_usb_device_controller/test_packet_inst/n129_s2  (
    .F(u_usb_device_controller_test_packet_inst_n129),
    .I0(u_usb_device_controller_test_packet_inst_cnt[8]),
    .I1(u_usb_device_controller_test_packet_inst_n129_6),
    .I2(u_usb_device_controller_test_packet_inst_cnt[9]),
    .I3(u_usb_device_controller_test_packet_inst_n127_7) 
);
defparam \u_usb_device_controller/test_packet_inst/n129_s2 .INIT=16'h7800;
  LUT3 \u_usb_device_controller/test_packet_inst/n130_s2  (
    .F(u_usb_device_controller_test_packet_inst_n130),
    .I0(u_usb_device_controller_test_packet_inst_n130_6),
    .I1(u_usb_device_controller_test_packet_inst_cnt[8]),
    .I2(u_usb_device_controller_test_packet_inst_n129_6) 
);
defparam \u_usb_device_controller/test_packet_inst/n130_s2 .INIT=8'h14;
  LUT4 \u_usb_device_controller/test_packet_inst/n131_s2  (
    .F(u_usb_device_controller_test_packet_inst_n131),
    .I0(u_usb_device_controller_test_packet_inst_cnt[6]),
    .I1(u_usb_device_controller_test_packet_inst_n131_8),
    .I2(u_usb_device_controller_test_packet_inst_n130_6),
    .I3(u_usb_device_controller_test_packet_inst_cnt[7]) 
);
defparam \u_usb_device_controller/test_packet_inst/n131_s2 .INIT=16'h0708;
  LUT3 \u_usb_device_controller/test_packet_inst/n132_s2  (
    .F(u_usb_device_controller_test_packet_inst_n132),
    .I0(u_usb_device_controller_test_packet_inst_n130_6),
    .I1(u_usb_device_controller_test_packet_inst_cnt[6]),
    .I2(u_usb_device_controller_test_packet_inst_n131_8) 
);
defparam \u_usb_device_controller/test_packet_inst/n132_s2 .INIT=8'h14;
  LUT4 \u_usb_device_controller/test_packet_inst/n133_s2  (
    .F(u_usb_device_controller_test_packet_inst_n133),
    .I0(u_usb_device_controller_test_packet_inst_n133_6),
    .I1(u_usb_device_controller_test_packet_inst_n133_7),
    .I2(u_usb_device_controller_test_packet_inst_n130_6),
    .I3(u_usb_device_controller_test_packet_inst_cnt[5]) 
);
defparam \u_usb_device_controller/test_packet_inst/n133_s2 .INIT=16'h0708;
  LUT4 \u_usb_device_controller/test_packet_inst/n134_s2  (
    .F(u_usb_device_controller_test_packet_inst_n134),
    .I0(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I1(u_usb_device_controller_test_packet_inst_n133_6),
    .I2(u_usb_device_controller_test_packet_inst_n130_6),
    .I3(u_usb_device_controller_test_packet_inst_cnt[4]) 
);
defparam \u_usb_device_controller/test_packet_inst/n134_s2 .INIT=16'h0708;
  LUT3 \u_usb_device_controller/test_packet_inst/n135_s2  (
    .F(u_usb_device_controller_test_packet_inst_n135),
    .I0(u_usb_device_controller_test_packet_inst_n130_6),
    .I1(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I2(u_usb_device_controller_test_packet_inst_n133_6) 
);
defparam \u_usb_device_controller/test_packet_inst/n135_s2 .INIT=8'h14;
  LUT4 \u_usb_device_controller/test_packet_inst/n136_s2  (
    .F(u_usb_device_controller_test_packet_inst_n136),
    .I0(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I2(u_usb_device_controller_test_packet_inst_n130_6),
    .I3(u_usb_device_controller_test_packet_inst_cnt[2]) 
);
defparam \u_usb_device_controller/test_packet_inst/n136_s2 .INIT=16'h0708;
  LUT3 \u_usb_device_controller/test_packet_inst/n137_s2  (
    .F(u_usb_device_controller_test_packet_inst_n137),
    .I0(u_usb_device_controller_test_packet_inst_n130_6),
    .I1(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[1]) 
);
defparam \u_usb_device_controller/test_packet_inst/n137_s2 .INIT=8'h14;
  LUT2 \u_usb_device_controller/test_packet_inst/n138_s2  (
    .F(u_usb_device_controller_test_packet_inst_n138),
    .I0(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I1(u_usb_device_controller_test_packet_inst_n130_6) 
);
defparam \u_usb_device_controller/test_packet_inst/n138_s2 .INIT=4'h1;
  LUT3 \u_usb_device_controller/test_packet_inst/n378_s0  (
    .F(u_usb_device_controller_test_packet_inst_n378),
    .I0(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dect),
    .I2(u_usb_device_controller_test_packet_inst_n378_4) 
);
defparam \u_usb_device_controller/test_packet_inst/n378_s0 .INIT=8'h40;
  LUT3 \u_usb_device_controller/u_usb_packet/n778_s0  (
    .F(u_usb_device_controller_u_usb_packet_n778),
    .I0(u_usb_device_controller_u_usb_packet_n640),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[7]),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n778_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/u_usb_packet/n779_s0  (
    .F(u_usb_device_controller_u_usb_packet_n779),
    .I0(u_usb_device_controller_u_usb_packet_n642),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[6]),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n779_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/u_usb_packet/n780_s0  (
    .F(u_usb_device_controller_u_usb_packet_n780),
    .I0(u_usb_device_controller_u_usb_packet_n644),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[5]),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n780_s0 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/u_usb_packet/n781_s0  (
    .F(u_usb_device_controller_u_usb_packet_n781),
    .I0(u_usb_device_controller_u_usb_packet_n646),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[4]),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n781_s0 .INIT=8'hAC;
  LUT4 \u_usb_device_controller/u_usb_packet/n782_s0  (
    .F(u_usb_device_controller_u_usb_packet_n782),
    .I0(u_usb_device_controller_u_usb_packet_n782_4),
    .I1(u_usb_device_controller_u_usb_packet_n782_5),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout[3]),
    .I3(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n782_s0 .INIT=16'h75F0;
  LUT3 \u_usb_device_controller/u_usb_packet/n783_s0  (
    .F(u_usb_device_controller_u_usb_packet_n783),
    .I0(u_usb_device_controller_u_usb_packet_n650),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[2]),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n783_s0 .INIT=8'hAC;
  LUT4 \u_usb_device_controller/u_usb_packet/n784_s0  (
    .F(u_usb_device_controller_u_usb_packet_n784),
    .I0(u_usb_device_controller_u_usb_packet_n784_4),
    .I1(u_usb_device_controller_u_usb_packet_n784_18),
    .I2(u_usb_device_controller_u_usb_packet_n784_6),
    .I3(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s0 .INIT=16'hD5F0;
  LUT4 \u_usb_device_controller/u_usb_packet/n785_s0  (
    .F(u_usb_device_controller_u_usb_packet_n785),
    .I0(u_usb_device_controller_u_usb_packet_n785_4),
    .I1(u_usb_device_controller_u_usb_packet_n784_18),
    .I2(u_usb_device_controller_u_usb_packet_n785_5),
    .I3(u_usb_device_controller_u_usb_packet_s_dataout_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n785_s0 .INIT=16'hD5F0;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s0  (
    .F(u_usb_device_controller_u_usb_packet_n912),
    .I0(u_usb_device_controller_u_usb_packet_n912_4),
    .I1(u_usb_device_controller_u_usb_packet_n912_5),
    .I2(u_usb_device_controller_u_usb_packet_n912_6),
    .I3(u_usb_device_controller_u_usb_packet_n912_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s0 .INIT=16'hFF80;
  LUT3 \u_usb_device_controller/u_usb_packet/n919_s0  (
    .F(u_usb_device_controller_u_usb_packet_n919),
    .I0(u_usb_device_controller_u_usb_packet_n784_20),
    .I1(u_usb_device_controller_u_usb_packet_n784_18),
    .I2(utmi_txready_i_d) 
);
defparam \u_usb_device_controller/u_usb_packet/n919_s0 .INIT=8'hF4;
  LUT3 \u_usb_device_controller/u_usb_packet/n920_s0  (
    .F(u_usb_device_controller_u_usb_packet_n920),
    .I0(u_usb_device_controller_u_usb_packet_n1454),
    .I1(u_usb_device_controller_u_usb_packet_n920_4),
    .I2(u_usb_device_controller_u_usb_packet_n920_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n920_s0 .INIT=8'hF1;
  LUT2 \u_usb_device_controller/usb_transact_inst/T_PING_s1  (
    .F(u_usb_device_controller_usb_transact_inst_T_PING),
    .I0(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I1(u_usb_device_controller_usb_transact_inst_s_ping) 
);
defparam \u_usb_device_controller/usb_transact_inst/T_PING_s1 .INIT=4'h4;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1041_s0  (
    .F(u_usb_device_controller_usb_transact_inst_n1041),
    .I0(u_usb_device_controller_usb_transact_inst_n1041_4),
    .I1(u_usb_device_controller_usb_transact_inst_n1041_8),
    .I2(u_usb_device_controller_usb_transact_inst_n1041_6) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1041_s0 .INIT=8'h80;
  LUT3 \u_usb_device_controller/usb_control_inst/n1629_s0  (
    .F(u_usb_device_controller_usb_control_inst_n1629),
    .I0(u_usb_device_controller_usb_control_inst_n1629_4),
    .I1(u_usb_device_controller_usb_control_inst_n1629_5),
    .I2(u_usb_device_controller_usb_control_inst_n1629_6) 
);
defparam \u_usb_device_controller/usb_control_inst/n1629_s0 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_control_inst/n2896_s0  (
    .F(u_usb_device_controller_usb_control_inst_n2896),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]),
    .I2(u_usb_device_controller_usb_control_inst_n2896_4),
    .I3(u_usb_device_controller_usb_control_inst_n2896_5) 
);
defparam \u_usb_device_controller/usb_control_inst/n2896_s0 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s19  (
    .F(u_usb_device_controller_u_usb_init_n212),
    .I0(u_usb_device_controller_u_usb_init_n212_28),
    .I1(u_usb_device_controller_u_usb_init_n212_29),
    .I2(u_usb_device_controller_u_usb_init_n212_61),
    .I3(u_usb_device_controller_u_usb_init_n212_31) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s19 .INIT=16'h88F0;
  LUT4 \u_usb_device_controller/u_usb_init/n215_s43  (
    .F(u_usb_device_controller_u_usb_init_n215),
    .I0(u_usb_device_controller_u_usb_init_n215_71),
    .I1(u_usb_device_controller_u_usb_init_s_state[2]),
    .I2(u_usb_device_controller_u_usb_init_s_state[3]),
    .I3(u_usb_device_controller_u_usb_init_n215_52) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s43 .INIT=16'h00EF;
  LUT4 \u_usb_device_controller/u_usb_init/n216_s42  (
    .F(u_usb_device_controller_u_usb_init_n216),
    .I0(u_usb_device_controller_u_usb_init_n216_49),
    .I1(u_usb_device_controller_u_usb_init_n414_4),
    .I2(u_usb_device_controller_u_usb_init_n216_56),
    .I3(u_usb_device_controller_u_usb_init_n216_51) 
);
defparam \u_usb_device_controller/u_usb_init/n216_s42 .INIT=16'hFFB0;
  LUT4 \u_usb_device_controller/usb_control_inst/n435_s11  (
    .F(u_usb_device_controller_usb_control_inst_n435),
    .I0(u_usb_device_controller_usb_control_inst_n435_16),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n435_17) 
);
defparam \u_usb_device_controller/usb_control_inst/n435_s11 .INIT=16'hF444;
  LUT4 \u_usb_device_controller/usb_control_inst/n436_s11  (
    .F(u_usb_device_controller_usb_control_inst_n436),
    .I0(u_usb_device_controller_usb_control_inst_n435_16),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[6]),
    .I3(u_usb_device_controller_usb_control_inst_n435_17) 
);
defparam \u_usb_device_controller/usb_control_inst/n436_s11 .INIT=16'hF444;
  LUT4 \u_usb_device_controller/usb_control_inst/n437_s11  (
    .F(u_usb_device_controller_usb_control_inst_n437),
    .I0(u_usb_device_controller_usb_control_inst_n435_16),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[5]),
    .I3(u_usb_device_controller_usb_control_inst_n435_17) 
);
defparam \u_usb_device_controller/usb_control_inst/n437_s11 .INIT=16'hF444;
  LUT4 \u_usb_device_controller/usb_control_inst/n438_s11  (
    .F(u_usb_device_controller_usb_control_inst_n438),
    .I0(u_usb_device_controller_usb_control_inst_n435_16),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[4]),
    .I3(u_usb_device_controller_usb_control_inst_n435_17) 
);
defparam \u_usb_device_controller/usb_control_inst/n438_s11 .INIT=16'hF444;
  LUT4 \u_usb_device_controller/usb_control_inst/n439_s11  (
    .F(u_usb_device_controller_usb_control_inst_n439),
    .I0(u_usb_device_controller_usb_control_inst_n435_16),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I3(u_usb_device_controller_usb_control_inst_n435_17) 
);
defparam \u_usb_device_controller/usb_control_inst/n439_s11 .INIT=16'hF444;
  LUT4 \u_usb_device_controller/usb_control_inst/n440_s11  (
    .F(u_usb_device_controller_usb_control_inst_n440),
    .I0(u_usb_device_controller_usb_control_inst_n435_16),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_n435_17) 
);
defparam \u_usb_device_controller/usb_control_inst/n440_s11 .INIT=16'hF444;
  LUT4 \u_usb_device_controller/usb_control_inst/n441_s11  (
    .F(u_usb_device_controller_usb_control_inst_n441),
    .I0(u_usb_device_controller_usb_control_inst_n435_16),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I3(u_usb_device_controller_usb_control_inst_n435_17) 
);
defparam \u_usb_device_controller/usb_control_inst/n441_s11 .INIT=16'hF444;
  LUT4 \u_usb_device_controller/usb_control_inst/n442_s11  (
    .F(u_usb_device_controller_usb_control_inst_n442),
    .I0(u_usb_device_controller_usb_control_inst_n435_16),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I3(u_usb_device_controller_usb_control_inst_n435_17) 
);
defparam \u_usb_device_controller/usb_control_inst/n442_s11 .INIT=16'hF444;
  LUT2 \u_usb_device_controller/u_usb_init/phy_linestate_rst_s1  (
    .F(u_usb_device_controller_u_usb_init_phy_linestate_rst),
    .I0(utmi_linestate_i_d[1]),
    .I1(utmi_linestate_i_d[0]) 
);
defparam \u_usb_device_controller/u_usb_init/phy_linestate_rst_s1 .INIT=4'hB;
  LUT2 \u_usb_device_controller/u_usb_packet/n328_s5  (
    .F(u_usb_device_controller_u_usb_packet_n328),
    .I0(u_usb_device_controller_u_usb_packet_n328_10),
    .I1(u_usb_device_controller_u_usb_packet_n328_11) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s5 .INIT=4'h8;
  LUT4 \u_usb_device_controller/usb_control_inst/n1836_s2  (
    .F(u_usb_device_controller_usb_control_inst_n1836),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I1(u_usb_device_controller_usb_control_inst_n1836_15),
    .I2(u_usb_device_controller_usb_control_inst_n1836_13),
    .I3(u_usb_device_controller_usb_control_inst_n1836_8) 
);
defparam \u_usb_device_controller/usb_control_inst/n1836_s2 .INIT=16'h8000;
  LUT3 \u_usb_device_controller/usb_control_inst/n1837_s2  (
    .F(u_usb_device_controller_usb_control_inst_n1837),
    .I0(u_usb_device_controller_usb_control_inst_n1836_15),
    .I1(u_usb_device_controller_usb_control_inst_n1837_6),
    .I2(u_usb_device_controller_usb_control_inst_n1837_7) 
);
defparam \u_usb_device_controller/usb_control_inst/n1837_s2 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_control_inst/n1864_s2  (
    .F(u_usb_device_controller_usb_control_inst_n1864),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I1(u_usb_device_controller_usb_control_inst_n1864_8),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .I3(u_usb_device_controller_usb_control_inst_n1699) 
);
defparam \u_usb_device_controller/usb_control_inst/n1864_s2 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/n2070_s2  (
    .F(u_usb_device_controller_usb_control_inst_n2070),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I3(u_usb_device_controller_usb_control_inst_n2067_6) 
);
defparam \u_usb_device_controller/usb_control_inst/n2070_s2 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/usb_control_inst/n1876_s1  (
    .F(u_usb_device_controller_usb_control_inst_n1876),
    .I0(u_usb_device_controller_usb_control_inst_n1876_9),
    .I1(u_usb_device_controller_usb_control_inst_n1876_13),
    .I2(u_usb_device_controller_usb_control_inst_n1876_11) 
);
defparam \u_usb_device_controller/usb_control_inst/n1876_s1 .INIT=8'h80;
  LUT2 \u_usb_device_controller/u_usb_init/n242_s1  (
    .F(u_usb_device_controller_u_usb_init_n242),
    .I0(reset_i_d),
    .I1(u_usb_device_controller_u_usb_init_v_clrtimer1) 
);
defparam \u_usb_device_controller/u_usb_init/n242_s1 .INIT=4'h4;
  LUT2 \u_usb_device_controller/u_usb_init/n280_s1  (
    .F(u_usb_device_controller_u_usb_init_n280),
    .I0(reset_i_d),
    .I1(u_usb_device_controller_u_usb_init_v_clrtimer2) 
);
defparam \u_usb_device_controller/u_usb_init/n280_s1 .INIT=4'h4;
  LUT2 \u_usb_device_controller/u_usb_packet/n800_s2  (
    .F(u_usb_device_controller_u_usb_packet_n800),
    .I0(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I1(u_usb_device_controller_u_usb_packet_n800_6) 
);
defparam \u_usb_device_controller/u_usb_packet/n800_s2 .INIT=4'hB;
  LUT4 \u_usb_device_controller/rxdat_d0_7_s3  (
    .F(u_usb_device_controller_rxdat_d0_7),
    .I0(u_usb_device_controller_rxdat_d0_7_9),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_n2393),
    .I3(u_usb_device_controller_rxdat_d0_7_10) 
);
defparam \u_usb_device_controller/rxdat_d0_7_s3 .INIT=16'hFFF4;
  LUT2 \u_usb_device_controller/u_usb_init/s_state_3_s3  (
    .F(u_usb_device_controller_u_usb_init_s_state_0),
    .I0(u_usb_device_controller_u_usb_init_s_state_3),
    .I1(u_usb_device_controller_u_usb_init_s_state_3_10) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s3 .INIT=4'h8;
  LUT3 \u_usb_device_controller/u_usb_packet/crc16_buf_15_s3  (
    .F(u_usb_device_controller_u_usb_packet_crc16_buf_15),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf_15_12),
    .I1(u_usb_device_controller_u_usb_packet_n784_18),
    .I2(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_15_s3 .INIT=8'h0D;
  LUT4 \u_usb_device_controller/usb_control_inst/s_answerlen_7_s2  (
    .F(u_usb_device_controller_usb_control_inst_s_answerlen_7),
    .I0(u_usb_device_controller_usb_control_inst_s_answerlen_7_7),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I2(u_usb_device_controller_usb_control_inst_n2067_6),
    .I3(u_usb_device_controller_usb_control_inst_s_setupptr[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerlen_7_s2 .INIT=16'h4000;
  LUT2 \u_usb_device_controller/n1619_s5  (
    .F(u_usb_device_controller_n1619),
    .I0(u_usb_device_controller_n384_10),
    .I1(u_usb_device_controller_n1585) 
);
defparam \u_usb_device_controller/n1619_s5 .INIT=4'hE;
  LUT2 \u_usb_device_controller/u_usb_packet/n615_s36  (
    .F(u_usb_device_controller_u_usb_packet_n615),
    .I0(u_usb_device_controller_u_usb_packet_n615_49),
    .I1(u_usb_device_controller_u_usb_packet_n615_42) 
);
defparam \u_usb_device_controller/u_usb_packet/n615_s36 .INIT=4'hB;
  LUT4 \u_usb_device_controller/u_usb_packet/s_dataout_7_s4  (
    .F(u_usb_device_controller_u_usb_packet_s_dataout_7),
    .I0(u_usb_device_controller_u_usb_packet_s_state[8]),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout_7_9),
    .I2(u_usb_device_controller_u_usb_packet_n615_49),
    .I3(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/s_dataout_7_s4 .INIT=16'h00F4;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1080_s40  (
    .F(u_usb_device_controller_usb_transact_inst_n1091),
    .I0(u_usb_device_controller_usb_transact_inst_n1080),
    .I1(u_usb_device_controller_usb_transact_inst_n1138_41),
    .I2(u_usb_device_controller_usb_transact_inst_n1080_46),
    .I3(u_usb_device_controller_usb_transact_inst_n1080_55) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1080_s40 .INIT=16'hEFFF;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1074_s15  (
    .F(u_usb_device_controller_usb_transact_inst_n1074_19),
    .I0(u_usb_device_controller_usb_transact_inst_n1074_22),
    .I1(u_usb_device_controller_usb_transact_inst_n1064_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1074_s15 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1072_s10  (
    .F(u_usb_device_controller_usb_transact_inst_n1072_15),
    .I0(u_usb_device_controller_usb_transact_inst_n1072_18),
    .I1(u_usb_device_controller_usb_transact_inst_n1072_19) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1072_s10 .INIT=4'hE;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1157_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I0(u_usb_device_controller_usb_transact_inst_n1157_26),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_27),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_28),
    .I3(u_usb_device_controller_usb_transact_inst_n1157_29) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1157_s18 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1670_s34  (
    .F(u_usb_device_controller_usb_control_inst_n1670),
    .I0(u_usb_device_controller_usb_control_inst_n1670_39),
    .I1(u_usb_device_controller_usb_control_inst_n1670_40),
    .I2(u_usb_device_controller_usb_control_inst_n1670_41),
    .I3(u_usb_device_controller_usb_control_inst_n1670_45) 
);
defparam \u_usb_device_controller/usb_control_inst/n1670_s34 .INIT=16'hBFFF;
  LUT4 \u_usb_device_controller/usb_control_inst/s_answerptr_7_s5  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_7_8),
    .I0(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerptr_7_11),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_12),
    .I3(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_7_s5 .INIT=16'h00F4;
  LUT4 \u_usb_device_controller/usb_control_inst/s_answerptr_5_s6  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_5),
    .I0(u_usb_device_controller_usb_control_inst_s_answerptr_5_10),
    .I1(u_usb_device_controller_usb_control_inst_s_answerptr_5_14),
    .I2(u_usb_device_controller_usb_control_inst_n1670_45),
    .I3(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_5_s6 .INIT=16'h00EF;
  LUT3 \u_usb_device_controller/u_usb_packet/s_state_11_s14  (
    .F(u_usb_device_controller_u_usb_packet_s_state_3),
    .I0(u_usb_device_controller_u_usb_packet_n800_6),
    .I1(u_usb_device_controller_u_usb_packet_n328_10),
    .I2(u_usb_device_controller_u_usb_packet_s_state_11) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_11_s14 .INIT=8'hD0;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_sof_s6  (
    .F(u_usb_device_controller_usb_transact_inst_s_sof_11),
    .I0(u_usb_device_controller_usb_transact_inst_s_sof_valid),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I2(u_usb_device_controller_usb_transact_inst_n1080_55),
    .I3(u_usb_device_controller_usb_transact_inst_n1111) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sof_s6 .INIT=16'hFF0B;
  LUT3 \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s4  (
    .F(u_usb_device_controller_usb_transact_inst_s_sendpid_0),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid_3_11),
    .I2(u_usb_device_controller_usb_transact_inst_s_sendpid_3_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s4 .INIT=8'h0B;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_1_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_1),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1701) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_1_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_2_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_2),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1703) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_2_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_3_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_3),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1705) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_3_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_4_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_4),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1707) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_4_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_5_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_5),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1709) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_5_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_6_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_6),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1711) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_6_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_7_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_7),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1713) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_7_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_8_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_8),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1715) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_8_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_9_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_9),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1717) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_9_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_10_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_10),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1719) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_10_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_11_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_11),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1721) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_11_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_12_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_12),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1723) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_12_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_13_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_13),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1725) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_13_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_14_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_14),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1727) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_14_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLRIN_15_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_15),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1729) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_15_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_1_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_1),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1731) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_1_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_2_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_2),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1733) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_2_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_3_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_3),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1735) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_3_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_4_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_4),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1737) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_4_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_5_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_5),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1739) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_5_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_6_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_6),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1741) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_6_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_7_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_7),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1743) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_7_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_8_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_8),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1745) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_8_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_9_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_9),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1747) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_9_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_10_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_10),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1749) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_10_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_11_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_11),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1751) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_11_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_12_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_12),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1753) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_12_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_13_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_13),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1755) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_13_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_14_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_14),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1757) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_14_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_CLROUT_15_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_CLROUT_15),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1759) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLROUT_15_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_1_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_1),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1761) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_1_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_2_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_2),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1763) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_2_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_3_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_3),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1765) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_3_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_4_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_4),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1767) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_4_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_5_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_5),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1769) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_5_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_6_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_6),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1771) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_6_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_7_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_7),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1773) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_7_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_8_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_8),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1775) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_8_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_9_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_9),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1777) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_9_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_10_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_10),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1779) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_10_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_11_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_11),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1781) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_11_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_12_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_12),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1783) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_12_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_13_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_13),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1785) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_13_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_14_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_14),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1787) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_14_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTIN_15_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTIN_15),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1789) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTIN_15_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_1_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_1),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1791) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_1_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_2_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_2),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1793) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_2_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_3_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_3),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1795) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_3_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_4_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_4),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1797) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_4_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_5_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_5),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1799) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_5_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_6_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_6),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1801) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_6_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_7_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_7),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1803) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_7_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_8_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_8),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1805) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_8_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_9_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_9),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1807) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_9_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_10_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_10),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1809) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_10_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_11_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_11),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1811) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_11_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_12_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_12),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1813) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_12_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_13_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_13),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1815) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_13_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_14_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_14),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1817) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_14_s4 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/C_SHLTOUT_15_s4  (
    .F(u_usb_device_controller_usb_control_inst_C_SHLTOUT_15),
    .I0(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I1(u_usb_device_controller_usb_control_inst_n1819) 
);
defparam \u_usb_device_controller/usb_control_inst/C_SHLTOUT_15_s4 .INIT=4'hE;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1068_s5  (
    .F(u_usb_device_controller_usb_transact_inst_n1068),
    .I0(u_usb_device_controller_usb_transact_inst_n1068_10),
    .I1(u_usb_device_controller_usb_transact_inst_n1068_16),
    .I2(u_usb_device_controller_usb_transact_inst_s_setup_2),
    .I3(u_usb_device_controller_usb_transact_inst_n1064_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1068_s5 .INIT=16'hBAF0;
  LUT4 \u_usb_device_controller/u_usb_packet/n640_s12  (
    .F(u_usb_device_controller_u_usb_packet_n640),
    .I0(u_usb_device_controller_u_usb_packet_n782_5),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[7]),
    .I2(u_usb_device_controller_u_usb_packet_n640_18),
    .I3(u_usb_device_controller_u_usb_packet_n640_19) 
);
defparam \u_usb_device_controller/u_usb_packet/n640_s12 .INIT=16'hF4FF;
  LUT3 \u_usb_device_controller/u_usb_packet/n642_s12  (
    .F(u_usb_device_controller_u_usb_packet_n642),
    .I0(u_usb_device_controller_u_usb_packet_n642_18),
    .I1(u_usb_device_controller_u_usb_packet_n642_19),
    .I2(u_usb_device_controller_u_usb_packet_n642_20) 
);
defparam \u_usb_device_controller/u_usb_packet/n642_s12 .INIT=8'h1F;
  LUT3 \u_usb_device_controller/u_usb_packet/n644_s12  (
    .F(u_usb_device_controller_u_usb_packet_n644),
    .I0(u_usb_device_controller_u_usb_packet_n644_18),
    .I1(u_usb_device_controller_u_usb_packet_n644_19),
    .I2(u_usb_device_controller_u_usb_packet_n644_20) 
);
defparam \u_usb_device_controller/u_usb_packet/n644_s12 .INIT=8'h1F;
  LUT4 \u_usb_device_controller/u_usb_packet/n646_s12  (
    .F(u_usb_device_controller_u_usb_packet_n646),
    .I0(u_usb_device_controller_u_usb_packet_n782_5),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[4]),
    .I2(u_usb_device_controller_u_usb_packet_n646_18),
    .I3(u_usb_device_controller_u_usb_packet_n646_19) 
);
defparam \u_usb_device_controller/u_usb_packet/n646_s12 .INIT=16'hF4FF;
  LUT4 \u_usb_device_controller/u_usb_packet/n650_s12  (
    .F(u_usb_device_controller_u_usb_packet_n650),
    .I0(u_usb_device_controller_u_usb_packet_n782_5),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[2]),
    .I2(u_usb_device_controller_u_usb_packet_n650_18),
    .I3(u_usb_device_controller_u_usb_packet_n650_19) 
);
defparam \u_usb_device_controller/u_usb_packet/n650_s12 .INIT=16'hF4FF;
  LUT4 \u_usb_device_controller/u_usb_packet/n652_s12  (
    .F(u_usb_device_controller_u_usb_packet_n652),
    .I0(u_usb_device_controller_u_usb_packet_n328_10),
    .I1(u_usb_device_controller_u_usb_packet_n626),
    .I2(u_usb_device_controller_u_usb_packet_n652_18),
    .I3(u_usb_device_controller_u_usb_packet_n784_4) 
);
defparam \u_usb_device_controller/u_usb_packet/n652_s12 .INIT=16'hF8FF;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1064_s10  (
    .F(u_usb_device_controller_usb_transact_inst_n1064),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I1(u_usb_device_controller_usb_transact_inst_n1064_18),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I3(u_usb_device_controller_usb_transact_inst_n1064_25) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1064_s10 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1066_s9  (
    .F(u_usb_device_controller_usb_transact_inst_n1066),
    .I0(u_usb_device_controller_usb_transact_inst_n1066_14),
    .I1(u_usb_device_controller_usb_transact_inst_n1064_18),
    .I2(u_usb_device_controller_usb_transact_inst_n1068_16),
    .I3(u_usb_device_controller_usb_transact_inst_s_out) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1066_s9 .INIT=16'h8F88;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1074_s16  (
    .F(u_usb_device_controller_usb_transact_inst_n1074),
    .I0(u_usb_device_controller_usb_transact_inst_n1068_16),
    .I1(u_usb_device_controller_usb_transact_inst_n1074_23),
    .I2(u_usb_device_controller_usb_transact_inst_n1074_24),
    .I3(u_usb_device_controller_usb_transact_inst_n1074_22) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1074_s16 .INIT=16'h4F44;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1070_s9  (
    .F(u_usb_device_controller_usb_transact_inst_n1070),
    .I0(u_usb_device_controller_usb_transact_inst_n1070_14),
    .I1(u_usb_device_controller_usb_transact_inst_n1070_18),
    .I2(u_usb_device_controller_usb_transact_inst_n1068_16),
    .I3(u_usb_device_controller_usb_transact_inst_s_ping) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1070_s9 .INIT=16'h4F44;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1163_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1163),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3_11),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I2(u_usb_device_controller_usb_transact_inst_n1163_24) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1163_s17 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_control_inst/n1672_s36  (
    .F(u_usb_device_controller_usb_control_inst_n1672),
    .I0(u_usb_device_controller_usb_control_inst_n1672_41),
    .I1(u_usb_device_controller_usb_control_inst_n1672_42),
    .I2(u_usb_device_controller_usb_control_inst_n1672_43),
    .I3(u_usb_device_controller_usb_control_inst_n1672_44) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s36 .INIT=16'h4F44;
  LUT4 \u_usb_device_controller/usb_control_inst/n1678_s34  (
    .F(u_usb_device_controller_usb_control_inst_n1678),
    .I0(u_usb_device_controller_usb_control_inst_n1678_46),
    .I1(u_usb_device_controller_usb_control_inst_n1678_40),
    .I2(u_usb_device_controller_usb_control_inst_n1678_41),
    .I3(u_usb_device_controller_usb_control_inst_n1672_44) 
);
defparam \u_usb_device_controller/usb_control_inst/n1678_s34 .INIT=16'hF400;
  LUT4 \u_usb_device_controller/usb_control_inst/n1680_s37  (
    .F(u_usb_device_controller_usb_control_inst_n1680),
    .I0(u_usb_device_controller_usb_control_inst_n1680_42),
    .I1(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I2(u_usb_device_controller_usb_control_inst_n1680_43),
    .I3(u_usb_device_controller_usb_control_inst_n1680_44) 
);
defparam \u_usb_device_controller/usb_control_inst/n1680_s37 .INIT=16'hFFF4;
  LUT4 \u_usb_device_controller/usb_control_inst/n1682_s34  (
    .F(u_usb_device_controller_usb_control_inst_n1682),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I1(u_usb_device_controller_usb_control_inst_n1682_39),
    .I2(u_usb_device_controller_usb_control_inst_n1629),
    .I3(u_usb_device_controller_usb_control_inst_n1682_40) 
);
defparam \u_usb_device_controller/usb_control_inst/n1682_s34 .INIT=16'h40FF;
  LUT4 \u_usb_device_controller/usb_control_inst/n1684_s34  (
    .F(u_usb_device_controller_usb_control_inst_n1684),
    .I0(u_usb_device_controller_usb_control_inst_n1682_39),
    .I1(u_usb_device_controller_usb_control_inst_n1684_39),
    .I2(u_usb_device_controller_usb_control_inst_n1836_15),
    .I3(u_usb_device_controller_usb_control_inst_n1684_40) 
);
defparam \u_usb_device_controller/usb_control_inst/n1684_s34 .INIT=16'hF888;
  LUT4 \u_usb_device_controller/usb_control_inst/n1686_s34  (
    .F(u_usb_device_controller_usb_control_inst_n1686),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I1(u_usb_device_controller_usb_control_inst_n1682_39),
    .I2(u_usb_device_controller_usb_control_inst_n1686_39),
    .I3(u_usb_device_controller_usb_control_inst_n1686_40) 
);
defparam \u_usb_device_controller/usb_control_inst/n1686_s34 .INIT=16'hFF40;
  LUT3 \u_usb_device_controller/usb_control_inst/n1688_s34  (
    .F(u_usb_device_controller_usb_control_inst_n1688),
    .I0(u_usb_device_controller_usb_control_inst_n1688_39),
    .I1(u_usb_device_controller_usb_control_inst_s_answerptr_7_12),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr_2_12) 
);
defparam \u_usb_device_controller/usb_control_inst/n1688_s34 .INIT=8'hF4;
  LUT4 \u_usb_device_controller/usb_control_inst/n1690_s29  (
    .F(u_usb_device_controller_usb_control_inst_n1690),
    .I0(u_usb_device_controller_usb_control_inst_n1690_34),
    .I1(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I2(u_usb_device_controller_usb_control_inst_n1690_35),
    .I3(u_usb_device_controller_usb_control_inst_n1690_36) 
);
defparam \u_usb_device_controller/usb_control_inst/n1690_s29 .INIT=16'hFFF4;
  LUT4 \u_usb_device_controller/usb_control_inst/n1701_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1701),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(u_usb_device_controller_usb_control_inst_n1701_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1701_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1703_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1703),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(u_usb_device_controller_usb_control_inst_n1701_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1703_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1705_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1705),
    .I0(u_usb_device_controller_usb_control_inst_n1701_17),
    .I1(u_usb_device_controller_usb_control_inst_n1705_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1705_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1707_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1707),
    .I0(u_usb_device_controller_usb_control_inst_n1701_17),
    .I1(u_usb_device_controller_usb_control_inst_n1707_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1707_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1709_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1709),
    .I0(u_usb_device_controller_usb_control_inst_n1701_17),
    .I1(u_usb_device_controller_usb_control_inst_n1709_19),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1709_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1711_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1711),
    .I0(u_usb_device_controller_usb_control_inst_n1701_17),
    .I1(u_usb_device_controller_usb_control_inst_n1711_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1711_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1713_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1713),
    .I0(u_usb_device_controller_usb_control_inst_n1701_17),
    .I1(u_usb_device_controller_usb_control_inst_n1713_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1713_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1715_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1715),
    .I0(u_usb_device_controller_usb_control_inst_n1715_16),
    .I1(u_usb_device_controller_usb_control_inst_n1715_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1715_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1717_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1717),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(u_usb_device_controller_usb_control_inst_n1715_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1717_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1719_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1719),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(u_usb_device_controller_usb_control_inst_n1715_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1719_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1721_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1721),
    .I0(u_usb_device_controller_usb_control_inst_n1705_16),
    .I1(u_usb_device_controller_usb_control_inst_n1715_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1721_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1723_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1723),
    .I0(u_usb_device_controller_usb_control_inst_n1707_16),
    .I1(u_usb_device_controller_usb_control_inst_n1715_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1723_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1725_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1725),
    .I0(u_usb_device_controller_usb_control_inst_n1709_19),
    .I1(u_usb_device_controller_usb_control_inst_n1715_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1725_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1727_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1727),
    .I0(u_usb_device_controller_usb_control_inst_n1711_16),
    .I1(u_usb_device_controller_usb_control_inst_n1715_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1727_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1729_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1729),
    .I0(u_usb_device_controller_usb_control_inst_n1713_16),
    .I1(u_usb_device_controller_usb_control_inst_n1715_17),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1729_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1731_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1731),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(u_usb_device_controller_usb_control_inst_n1731_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1731_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1733_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1733),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(u_usb_device_controller_usb_control_inst_n1731_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1733_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1735_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1735),
    .I0(u_usb_device_controller_usb_control_inst_n1705_16),
    .I1(u_usb_device_controller_usb_control_inst_n1731_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1735_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1737_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1737),
    .I0(u_usb_device_controller_usb_control_inst_n1707_16),
    .I1(u_usb_device_controller_usb_control_inst_n1731_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1737_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1739_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1739),
    .I0(u_usb_device_controller_usb_control_inst_n1709_19),
    .I1(u_usb_device_controller_usb_control_inst_n1731_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1739_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1741_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1741),
    .I0(u_usb_device_controller_usb_control_inst_n1711_16),
    .I1(u_usb_device_controller_usb_control_inst_n1731_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1741_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1743_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1743),
    .I0(u_usb_device_controller_usb_control_inst_n1713_16),
    .I1(u_usb_device_controller_usb_control_inst_n1731_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1743_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1745_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1745),
    .I0(u_usb_device_controller_usb_control_inst_n1715_16),
    .I1(u_usb_device_controller_usb_control_inst_n1745_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1745_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1747_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1747),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(u_usb_device_controller_usb_control_inst_n1745_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1747_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1749_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1749),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(u_usb_device_controller_usb_control_inst_n1745_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1749_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1751_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1751),
    .I0(u_usb_device_controller_usb_control_inst_n1705_16),
    .I1(u_usb_device_controller_usb_control_inst_n1745_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1751_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1753_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1753),
    .I0(u_usb_device_controller_usb_control_inst_n1707_16),
    .I1(u_usb_device_controller_usb_control_inst_n1745_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1753_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1755_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1755),
    .I0(u_usb_device_controller_usb_control_inst_n1709_19),
    .I1(u_usb_device_controller_usb_control_inst_n1745_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1755_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1757_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1757),
    .I0(u_usb_device_controller_usb_control_inst_n1711_16),
    .I1(u_usb_device_controller_usb_control_inst_n1745_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1757_s11 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1759_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1759),
    .I0(u_usb_device_controller_usb_control_inst_n1713_16),
    .I1(u_usb_device_controller_usb_control_inst_n1745_16),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1701_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1759_s11 .INIT=16'hF800;
  LUT3 \u_usb_device_controller/usb_control_inst/n1646_s6  (
    .F(u_usb_device_controller_usb_control_inst_n1646),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[6]),
    .I1(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I2(u_usb_device_controller_usb_control_inst_n1670_39) 
);
defparam \u_usb_device_controller/usb_control_inst/n1646_s6 .INIT=8'h60;
  LUT4 \u_usb_device_controller/usb_control_inst/n1649_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1649),
    .I0(u_usb_device_controller_usb_control_inst_n1649_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[5]),
    .I2(u_usb_device_controller_usb_control_inst_n1649_17),
    .I3(u_usb_device_controller_usb_control_inst_n1649_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1649_s11 .INIT=16'hBEAA;
  LUT4 \u_usb_device_controller/usb_control_inst/n1652_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1652),
    .I0(u_usb_device_controller_usb_control_inst_n1652_16),
    .I1(u_usb_device_controller_usb_control_inst_n1652_24),
    .I2(u_usb_device_controller_usb_control_inst_n1652_18),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscoff[4]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1652_s11 .INIT=16'hA30C;
  LUT4 \u_usb_device_controller/usb_control_inst/n1655_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1655),
    .I0(u_usb_device_controller_usb_control_inst_n1652_16),
    .I1(u_usb_device_controller_usb_control_inst_n1655_18),
    .I2(u_usb_device_controller_usb_control_inst_n1652_18),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscoff[3]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1655_s11 .INIT=16'hA30C;
  LUT4 \u_usb_device_controller/usb_control_inst/n1658_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1658),
    .I0(u_usb_device_controller_usb_control_inst_n1652_16),
    .I1(u_usb_device_controller_usb_control_inst_n1658_16),
    .I2(u_usb_device_controller_usb_control_inst_n1652_18),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscoff[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1658_s11 .INIT=16'hA30C;
  LUT4 \u_usb_device_controller/usb_control_inst/n1661_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1661),
    .I0(u_usb_device_controller_usb_control_inst_n1661_16),
    .I1(u_usb_device_controller_usb_control_inst_n1661_17),
    .I2(u_usb_device_controller_usb_control_inst_n1661_18),
    .I3(u_usb_device_controller_usb_control_inst_n1661_19) 
);
defparam \u_usb_device_controller/usb_control_inst/n1661_s11 .INIT=16'hFFF8;
  LUT3 \u_usb_device_controller/usb_control_inst/n1664_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1664),
    .I0(u_usb_device_controller_usb_control_inst_n1652_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I2(u_usb_device_controller_usb_control_inst_n1652_18) 
);
defparam \u_usb_device_controller/usb_control_inst/n1664_s11 .INIT=8'h83;
  LUT3 \u_usb_device_controller/usb_control_inst/n1696_s8  (
    .F(u_usb_device_controller_usb_control_inst_n1696),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .I2(u_usb_device_controller_usb_control_inst_n1836_15) 
);
defparam \u_usb_device_controller/usb_control_inst/n1696_s8 .INIT=8'h60;
  LUT3 \u_usb_device_controller/u_usb_packet/n626_s36  (
    .F(u_usb_device_controller_u_usb_packet_n626),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_u_usb_packet_n626_42),
    .I2(u_usb_device_controller_u_usb_packet_n626_48) 
);
defparam \u_usb_device_controller/u_usb_packet/n626_s36 .INIT=8'hD0;
  LUT3 \u_usb_device_controller/u_usb_packet/n628_s42  (
    .F(u_usb_device_controller_u_usb_packet_n628),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I2(u_usb_device_controller_u_usb_packet_n628_47) 
);
defparam \u_usb_device_controller/u_usb_packet/n628_s42 .INIT=8'h40;
  LUT3 \u_usb_device_controller/u_usb_packet/n630_s42  (
    .F(u_usb_device_controller_u_usb_packet_n630),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I2(u_usb_device_controller_u_usb_packet_n628_47) 
);
defparam \u_usb_device_controller/u_usb_packet/n630_s42 .INIT=8'h80;
  LUT2 \u_usb_device_controller/u_usb_packet/n632_s42  (
    .F(u_usb_device_controller_u_usb_packet_n632),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I1(u_usb_device_controller_u_usb_packet_n628_47) 
);
defparam \u_usb_device_controller/u_usb_packet/n632_s42 .INIT=4'h4;
  LUT4 \u_usb_device_controller/u_usb_packet/n633_s34  (
    .F(u_usb_device_controller_u_usb_packet_n633),
    .I0(u_usb_device_controller_u_usb_packet_n328_11),
    .I1(u_usb_device_controller_u_usb_packet_n800_6),
    .I2(u_usb_device_controller_u_usb_packet_n328_10),
    .I3(u_usb_device_controller_u_usb_packet_n633_39) 
);
defparam \u_usb_device_controller/u_usb_packet/n633_s34 .INIT=16'h40FF;
  LUT2 \u_usb_device_controller/u_usb_packet/n635_s36  (
    .F(u_usb_device_controller_u_usb_packet_n635),
    .I0(u_usb_device_controller_u_usb_init_usbp_chirpk),
    .I1(u_usb_device_controller_u_usb_packet_n784_18) 
);
defparam \u_usb_device_controller/u_usb_packet/n635_s36 .INIT=4'h8;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1086_s39  (
    .F(u_usb_device_controller_usb_transact_inst_n1086),
    .I0(u_usb_device_controller_usb_transact_inst_n1086_52),
    .I1(u_usb_device_controller_usb_transact_inst_n1086_48),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[12]),
    .I3(u_usb_device_controller_usb_transact_inst_n1086_50) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1086_s39 .INIT=16'hF888;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1088_s39  (
    .F(u_usb_device_controller_usb_transact_inst_n1088),
    .I0(u_usb_device_controller_usb_transact_inst_n1086_52),
    .I1(u_usb_device_controller_usb_transact_inst_n1088_44),
    .I2(u_usb_device_controller_usb_transact_inst_n1088_45),
    .I3(u_usb_device_controller_u_usb_packet_usbp_rxact) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1088_s39 .INIT=16'h8F88;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1090_s41  (
    .F(u_usb_device_controller_usb_transact_inst_n1090),
    .I0(u_usb_device_controller_usb_transact_inst_n1090_46),
    .I1(u_usb_device_controller_usb_transact_inst_n1064_16),
    .I2(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I3(u_usb_device_controller_usb_transact_inst_n1088_45) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1090_s41 .INIT=16'h444F;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1093_s46  (
    .F(u_usb_device_controller_usb_transact_inst_n1093),
    .I0(u_usb_device_controller_usb_transact_inst_n1093_51),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .I2(u_usb_device_controller_usb_transact_inst_n1163) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1093_s46 .INIT=8'hF4;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1095_s39  (
    .F(u_usb_device_controller_usb_transact_inst_n1095),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I1(u_usb_device_controller_usb_transact_inst_n1095_44),
    .I2(u_usb_device_controller_usb_transact_inst_n1095_45),
    .I3(u_usb_device_controller_usb_transact_inst_n1095_46) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1095_s39 .INIT=16'hF444;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1097_s42  (
    .F(u_usb_device_controller_usb_transact_inst_n1097),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[6]),
    .I1(u_usb_device_controller_usb_transact_inst_n1086_50),
    .I2(u_usb_device_controller_usb_transact_inst_n1565) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1097_s42 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1101_s39  (
    .F(u_usb_device_controller_usb_transact_inst_n1101),
    .I0(u_usb_device_controller_usb_transact_inst_n1095_46),
    .I1(u_usb_device_controller_usb_transact_inst_n1074_22),
    .I2(u_usb_device_controller_usb_transact_inst_n1101_44) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1101_s39 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1103_s40  (
    .F(u_usb_device_controller_usb_transact_inst_n1103),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[3]),
    .I1(u_usb_device_controller_usb_transact_inst_n1086_50),
    .I2(u_usb_device_controller_usb_transact_inst_s_endpt_3) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1103_s40 .INIT=8'hF8;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1105_s42  (
    .F(u_usb_device_controller_usb_transact_inst_n1105),
    .I0(u_usb_device_controller_usb_transact_inst_n1105_47),
    .I1(u_usb_device_controller_usb_transact_inst_s_endpt_0_9),
    .I2(u_usb_device_controller_usb_transact_inst_n1105_48),
    .I3(u_usb_device_controller_usb_transact_inst_n1041) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1105_s42 .INIT=16'hF444;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1107_s41  (
    .F(u_usb_device_controller_usb_transact_inst_n1107),
    .I0(u_usb_device_controller_usb_transact_inst_n1093_51),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[1]),
    .I2(u_usb_device_controller_usb_transact_inst_n1107_48) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1107_s41 .INIT=8'hF4;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1109_s42  (
    .F(u_usb_device_controller_usb_transact_inst_n1109),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I1(u_usb_device_controller_usb_transact_inst_n1138_24),
    .I2(u_usb_device_controller_usb_transact_inst_n1109_47),
    .I3(u_usb_device_controller_usb_transact_inst_n1109_48) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1109_s42 .INIT=16'hF8FF;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1138_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1138),
    .I0(u_usb_device_controller_usb_transact_inst_n1138_39),
    .I1(u_usb_device_controller_usb_transact_inst_n1138_43),
    .I2(u_usb_device_controller_usb_transact_inst_n1138_29),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_30) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s18 .INIT=16'hFFF8;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1142_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1142),
    .I0(u_usb_device_controller_usb_transact_inst_n1142_25),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[6]),
    .I2(u_usb_device_controller_usb_transact_inst_n1142_23),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_43) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1142_s17 .INIT=16'h7D55;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1144_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1144),
    .I0(u_usb_device_controller_usb_transact_inst_n1142_23),
    .I1(u_usb_device_controller_usb_transact_inst_n1138_43),
    .I2(u_usb_device_controller_usb_transact_inst_n1144_22),
    .I3(u_usb_device_controller_usb_transact_inst_n1142_25) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1144_s17 .INIT=16'hF8FF;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1146_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1146),
    .I0(u_usb_device_controller_usb_transact_inst_n1142_25),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[4]),
    .I2(u_usb_device_controller_usb_transact_inst_n1146_22),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_43) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1146_s17 .INIT=16'h7D55;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1148_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1148),
    .I0(u_usb_device_controller_usb_transact_inst_n1138_43),
    .I1(u_usb_device_controller_usb_transact_inst_n1146_22),
    .I2(u_usb_device_controller_usb_transact_inst_n1148_22),
    .I3(u_usb_device_controller_usb_transact_inst_n1148_25) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1148_s17 .INIT=16'hF8FF;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1150_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1150),
    .I0(u_usb_device_controller_usb_transact_inst_n1148_25),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[2]),
    .I2(u_usb_device_controller_usb_transact_inst_n1150_22),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_43) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1150_s17 .INIT=16'h7D55;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1152_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1152),
    .I0(u_usb_device_controller_usb_transact_inst_n1138_43),
    .I1(u_usb_device_controller_usb_transact_inst_n1150_22),
    .I2(u_usb_device_controller_usb_transact_inst_n1152_22),
    .I3(u_usb_device_controller_usb_transact_inst_n1148_25) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1152_s17 .INIT=16'hF8FF;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1154_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1154),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[0]),
    .I1(u_usb_device_controller_usb_transact_inst_n1138_43),
    .I2(u_usb_device_controller_usb_transact_inst_n1142_25) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1154_s17 .INIT=8'h4F;
  LUT4 \u_usb_device_controller/n1615_s9  (
    .F(u_usb_device_controller_n1615),
    .I0(u_usb_device_controller_n1585),
    .I1(u_usb_device_controller_usb_transact_inst_txpop_o_d),
    .I2(u_usb_device_controller_n1615_15),
    .I3(u_usb_device_controller_s_bufptr[0]) 
);
defparam \u_usb_device_controller/n1615_s9 .INIT=16'h30EA;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1076_s14  (
    .F(u_usb_device_controller_usb_transact_inst_n1076),
    .I0(u_usb_device_controller_usb_transact_inst_n1076_21),
    .I1(u_usb_device_controller_usb_transact_inst_n1074_22),
    .I2(u_usb_device_controller_usb_transact_inst_n1076_24) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1076_s14 .INIT=8'hF8;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1072_s11  (
    .F(u_usb_device_controller_usb_transact_inst_n1072),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I1(u_usb_device_controller_usb_transact_inst_n1095_46),
    .I2(u_usb_device_controller_usb_transact_inst_n1072_19),
    .I3(u_usb_device_controller_usb_transact_inst_n1072_20) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1072_s11 .INIT=16'hFFE0;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1157_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1157),
    .I0(u_usb_device_controller_usb_transact_inst_n1157_30),
    .I1(u_usb_device_controller_usb_transact_inst_n1163),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_31) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1157_s19 .INIT=8'hF4;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1159_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1159),
    .I0(u_usb_device_controller_usb_transact_inst_n1159_25),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid_3_23),
    .I2(u_usb_device_controller_usb_transact_inst_n1159_26) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1159_s19 .INIT=8'h01;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1161_s10  (
    .F(u_usb_device_controller_usb_transact_inst_n1161),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_0),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[1]),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1161_s10 .INIT=8'hE0;
  LUT4 \u_usb_device_controller/usb_control_inst/n1860_s23  (
    .F(u_usb_device_controller_usb_control_inst_n1860),
    .I0(u_usb_device_controller_usb_control_inst_n1860_29),
    .I1(u_usb_device_controller_usb_control_inst_n1876_13),
    .I2(u_usb_device_controller_usb_control_inst_n1864_8),
    .I3(u_usb_device_controller_usb_control_inst_n1860_30) 
);
defparam \u_usb_device_controller/usb_control_inst/n1860_s23 .INIT=16'hFF80;
  LUT3 \u_usb_device_controller/n1241_s61  (
    .F(u_usb_device_controller_n1241_60),
    .I0(u_usb_device_controller_halt_out[2]),
    .I1(u_usb_device_controller_halt_out[3]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1241_s61 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1242_s61  (
    .F(u_usb_device_controller_n1242_60),
    .I0(u_usb_device_controller_halt_in[2]),
    .I1(u_usb_device_controller_halt_in[3]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1242_s61 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1243_s61  (
    .F(u_usb_device_controller_n1243_60),
    .I0(u_usb_device_controller_osync[2]),
    .I1(u_usb_device_controller_osync[3]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1243_s61 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n1244_s61  (
    .F(u_usb_device_controller_n1244_60),
    .I0(u_usb_device_controller_isync[2]),
    .I1(u_usb_device_controller_isync[3]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]) 
);
defparam \u_usb_device_controller/n1244_s61 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n385_s2  (
    .F(u_usb_device_controller_n385_6),
    .I0(u_usb_device_controller_n385_7),
    .I1(u_usb_device_controller_n385_10),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n385_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n443_s2  (
    .F(u_usb_device_controller_n443_6),
    .I0(u_usb_device_controller_n443_7),
    .I1(u_usb_device_controller_n443_10),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n443_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n503_s2  (
    .F(u_usb_device_controller_n503_6),
    .I0(u_usb_device_controller_n503_7),
    .I1(u_usb_device_controller_n503_10),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n503_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n561_s2  (
    .F(u_usb_device_controller_n561_6),
    .I0(u_usb_device_controller_n561_7),
    .I1(u_usb_device_controller_n561_10),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n561_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n621_s2  (
    .F(u_usb_device_controller_n621_6),
    .I0(u_usb_device_controller_n385_7),
    .I1(u_usb_device_controller_n621_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n621_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n681_s2  (
    .F(u_usb_device_controller_n681_6),
    .I0(u_usb_device_controller_n443_7),
    .I1(u_usb_device_controller_n681_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n681_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n743_s2  (
    .F(u_usb_device_controller_n743_6),
    .I0(u_usb_device_controller_n503_7),
    .I1(u_usb_device_controller_n743_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n743_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n801_s2  (
    .F(u_usb_device_controller_n801_6),
    .I0(u_usb_device_controller_n561_7),
    .I1(u_usb_device_controller_n801_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n801_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n861_s2  (
    .F(u_usb_device_controller_n861_6),
    .I0(u_usb_device_controller_n385_7),
    .I1(u_usb_device_controller_n861_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n861_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n921_s2  (
    .F(u_usb_device_controller_n921_6),
    .I0(u_usb_device_controller_n443_7),
    .I1(u_usb_device_controller_n921_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n921_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n983_s2  (
    .F(u_usb_device_controller_n983_6),
    .I0(u_usb_device_controller_n503_7),
    .I1(u_usb_device_controller_n983_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n983_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n1043_s2  (
    .F(u_usb_device_controller_n1043_6),
    .I0(u_usb_device_controller_n561_7),
    .I1(u_usb_device_controller_n1043_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1043_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n1105_s2  (
    .F(u_usb_device_controller_n1105_6),
    .I0(u_usb_device_controller_n385_7),
    .I1(u_usb_device_controller_n1105_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1105_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n1167_s2  (
    .F(u_usb_device_controller_n1167_6),
    .I0(u_usb_device_controller_n443_7),
    .I1(u_usb_device_controller_n1167_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1167_s2 .INIT=8'hF8;
  LUT3 \u_usb_device_controller/n1231_s2  (
    .F(u_usb_device_controller_n1231_6),
    .I0(u_usb_device_controller_n503_7),
    .I1(u_usb_device_controller_n1231_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1231_s2 .INIT=8'hF8;
  LUT4 \u_usb_device_controller/test_packet_inst/cnt_11_s3  (
    .F(u_usb_device_controller_test_packet_inst_cnt_11),
    .I0(utmi_txready_i_d),
    .I1(u_usb_device_controller_test_packet_inst_cnt_11_9),
    .I2(u_usb_device_controller_test_packet_inst_cnt_11_10),
    .I3(u_usb_device_controller_test_packet_inst_test_en_dly_Z) 
);
defparam \u_usb_device_controller/test_packet_inst/cnt_11_s3 .INIT=16'hB0FF;
  LUT2 \u_usb_device_controller/test_packet_inst/test_data_6_s3  (
    .F(u_usb_device_controller_test_packet_inst_test_data_7),
    .I0(u_usb_device_controller_test_packet_inst_test_data_6),
    .I1(u_usb_device_controller_test_packet_inst_test_data_6_8) 
);
defparam \u_usb_device_controller/test_packet_inst/test_data_6_s3 .INIT=4'hB;
  LUT4 \u_usb_device_controller/test_packet_inst/test_data_val_s3  (
    .F(u_usb_device_controller_test_packet_inst_test_data_val),
    .I0(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I1(u_usb_device_controller_test_packet_inst_test_data_val_9),
    .I2(u_usb_device_controller_test_packet_inst_test_data_6_8),
    .I3(u_usb_device_controller_test_packet_inst_test_data_6) 
);
defparam \u_usb_device_controller/test_packet_inst/test_data_val_s3 .INIT=16'hFF07;
  LUT3 \u_usb_device_controller/u_usb_init/s_state_1_s8  (
    .F(u_usb_device_controller_u_usb_init_s_state_1),
    .I0(u_usb_device_controller_u_usb_init_s_state_3_10),
    .I1(u_usb_device_controller_u_usb_init_s_state[2]),
    .I2(u_usb_device_controller_u_usb_init_s_state_3) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_1_s8 .INIT=8'hB0;
  LUT2 \u_usb_device_controller/u_usb_init/n218_s22  (
    .F(u_usb_device_controller_u_usb_init_n218),
    .I0(u_usb_device_controller_u_usb_init_s_state[1]),
    .I1(u_usb_device_controller_u_usb_init_s_state[2]) 
);
defparam \u_usb_device_controller/u_usb_init/n218_s22 .INIT=4'h8;
  LUT2 \u_usb_device_controller/test_packet_inst/n319_s3  (
    .F(u_usb_device_controller_test_packet_inst_n319),
    .I0(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I1(u_usb_device_controller_test_packet_inst_cnt_11_9) 
);
defparam \u_usb_device_controller/test_packet_inst/n319_s3 .INIT=4'h8;
  LUT4 \u_usb_device_controller/test_packet_inst/n318_s3  (
    .F(u_usb_device_controller_test_packet_inst_n318),
    .I0(u_usb_device_controller_test_packet_inst_n318_8),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_test_packet_inst_n318_9),
    .I3(u_usb_device_controller_test_packet_inst_n318_10) 
);
defparam \u_usb_device_controller/test_packet_inst/n318_s3 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/test_packet_inst/n317_s4  (
    .F(u_usb_device_controller_test_packet_inst_n317),
    .I0(u_usb_device_controller_test_packet_inst_test_data_6),
    .I1(u_usb_device_controller_test_packet_inst_n317_9),
    .I2(u_usb_device_controller_test_packet_inst_n317_10),
    .I3(u_usb_device_controller_test_packet_inst_n318_10) 
);
defparam \u_usb_device_controller/test_packet_inst/n317_s4 .INIT=16'hFFE0;
  LUT4 \u_usb_device_controller/test_packet_inst/n312_s3  (
    .F(u_usb_device_controller_test_packet_inst_n312),
    .I0(u_usb_device_controller_test_packet_inst_n312_8),
    .I1(u_usb_device_controller_test_packet_inst_n312_9),
    .I2(u_usb_device_controller_test_packet_inst_n312_10),
    .I3(u_usb_device_controller_test_packet_inst_n318_10) 
);
defparam \u_usb_device_controller/test_packet_inst/n312_s3 .INIT=16'hFFB0;
  LUT3 \u_usb_device_controller/test_packet_inst/n311_s4  (
    .F(u_usb_device_controller_test_packet_inst_n311),
    .I0(u_usb_device_controller_test_packet_inst_n311_9),
    .I1(u_usb_device_controller_test_packet_inst_n317_10),
    .I2(u_usb_device_controller_test_packet_inst_n318_10) 
);
defparam \u_usb_device_controller/test_packet_inst/n311_s4 .INIT=8'hF4;
  LUT2 \u_usb_device_controller/n1244_s60  (
    .F(u_usb_device_controller_n1244_62),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_isync[1]) 
);
defparam \u_usb_device_controller/n1244_s60 .INIT=4'h8;
  LUT2 \u_usb_device_controller/n1243_s60  (
    .F(u_usb_device_controller_n1243_62),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_osync[1]) 
);
defparam \u_usb_device_controller/n1243_s60 .INIT=4'h8;
  LUT2 \u_usb_device_controller/n1242_s60  (
    .F(u_usb_device_controller_n1242_62),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_halt_in[1]) 
);
defparam \u_usb_device_controller/n1242_s60 .INIT=4'h8;
  LUT2 \u_usb_device_controller/n1241_s60  (
    .F(u_usb_device_controller_n1241_62),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_halt_out[1]) 
);
defparam \u_usb_device_controller/n1241_s60 .INIT=4'h8;
  LUT3 \u_usb_device_controller/u_usb_init/n208_s21  (
    .F(u_usb_device_controller_u_usb_init_n208),
    .I0(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I1(u_usb_device_controller_u_usb_init_s_state[1]),
    .I2(u_usb_device_controller_u_usb_init_n210) 
);
defparam \u_usb_device_controller/u_usb_init/n208_s21 .INIT=8'h07;
  LUT2 \u_usb_device_controller/u_usb_init/n222_s19  (
    .F(u_usb_device_controller_u_usb_init_n222),
    .I0(u_usb_device_controller_u_usb_init_s_chirpcnt[0]),
    .I1(u_usb_device_controller_u_usb_init_s_state[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n222_s19 .INIT=4'h4;
  LUT3 \u_usb_device_controller/u_usb_init/n221_s19  (
    .F(u_usb_device_controller_u_usb_init_n221),
    .I0(u_usb_device_controller_u_usb_init_s_chirpcnt[0]),
    .I1(u_usb_device_controller_u_usb_init_s_chirpcnt[1]),
    .I2(u_usb_device_controller_u_usb_init_s_state[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n221_s19 .INIT=8'h60;
  LUT4 \u_usb_device_controller/u_usb_init/n220_s19  (
    .F(u_usb_device_controller_u_usb_init_n220),
    .I0(u_usb_device_controller_u_usb_init_s_chirpcnt[0]),
    .I1(u_usb_device_controller_u_usb_init_s_chirpcnt[1]),
    .I2(u_usb_device_controller_u_usb_init_s_chirpcnt[2]),
    .I3(u_usb_device_controller_u_usb_init_s_state[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n220_s19 .INIT=16'h7800;
  LUT4 \u_usb_device_controller/u_usb_init/n213_s19  (
    .F(u_usb_device_controller_u_usb_init_n213),
    .I0(u_usb_device_controller_u_usb_init_s_state[2]),
    .I1(u_usb_device_controller_u_usb_init_n215_71),
    .I2(u_usb_device_controller_u_usb_init_s_state[3]),
    .I3(u_usb_device_controller_u_usb_init_n213_28) 
);
defparam \u_usb_device_controller/u_usb_init/n213_s19 .INIT=16'hFF40;
  LUT2 \u_usb_device_controller/u_usb_init/n219_s19  (
    .F(u_usb_device_controller_u_usb_init_n219),
    .I0(u_usb_device_controller_u_usb_init_s_state[3]),
    .I1(u_usb_device_controller_u_usb_init_n219_28) 
);
defparam \u_usb_device_controller/u_usb_init/n219_s19 .INIT=4'h4;
  LUT4 \u_usb_device_controller/n1534_s18  (
    .F(u_usb_device_controller_n1534),
    .I0(u_usb_device_controller_n1534_26),
    .I1(u_usb_device_controller_n1534_37),
    .I2(u_usb_device_controller_n1534_28),
    .I3(u_usb_device_controller_n1534_29) 
);
defparam \u_usb_device_controller/n1534_s18 .INIT=16'hFF0E;
  LUT4 \u_usb_device_controller/n1529_s17  (
    .F(u_usb_device_controller_n1529),
    .I0(u_usb_device_controller_n1529_24),
    .I1(u_usb_device_controller_n1529_25),
    .I2(u_usb_device_controller_n1529_26),
    .I3(u_usb_device_controller_n1529_31) 
);
defparam \u_usb_device_controller/n1529_s17 .INIT=16'hFFF8;
  LUT4 \u_usb_device_controller/n1524_s17  (
    .F(u_usb_device_controller_n1524),
    .I0(u_usb_device_controller_n1524_27),
    .I1(u_usb_device_controller_n1585_4),
    .I2(u_usb_device_controller_n1524_25),
    .I3(u_usb_device_controller_n1534_37) 
);
defparam \u_usb_device_controller/n1524_s17 .INIT=16'hFFF4;
  LUT4 \u_usb_device_controller/n1519_s20  (
    .F(u_usb_device_controller_n1519),
    .I0(u_usb_device_controller_usb_transact_inst_s_out_valid),
    .I1(u_usb_device_controller_cur_state[3]),
    .I2(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I3(u_usb_device_controller_n1519_32) 
);
defparam \u_usb_device_controller/n1519_s20 .INIT=16'h0D00;
  LUT2 \u_usb_device_controller/utmi_opmode_o_d_0_s  (
    .F(u_usb_device_controller_utmi_opmode_o_d[0]),
    .I0(u_usb_device_controller_u_usb_init_usbi_opmode[0]),
    .I1(u_usb_device_controller_utmi_txvalid_o_d_8) 
);
defparam \u_usb_device_controller/utmi_opmode_o_d_0_s .INIT=4'h8;
  LUT3 \u_usb_device_controller/usbc_dsclen_1_s8  (
    .F(u_usb_device_controller_usbc_dsclen_1),
    .I0(u_usb_device_controller_usbc_dsclen_0_28),
    .I1(u_usb_device_controller_usbc_dsclen_1_14),
    .I2(u_usb_device_controller_usbc_dsclen_1_15) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s8 .INIT=8'h01;
  LUT4 \u_usb_device_controller/usbc_dsclen_2_s8  (
    .F(u_usb_device_controller_usbc_dsclen_2),
    .I0(u_usb_device_controller_usbc_dsclen_2_14),
    .I1(u_usb_device_controller_usbc_dsclen_2_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_2_s8 .INIT=16'h0305;
  LUT2 \u_usb_device_controller/usbc_dsclen_3_s8  (
    .F(u_usb_device_controller_usbc_dsclen_3),
    .I0(u_usb_device_controller_usbc_dsclen_0_28),
    .I1(u_usb_device_controller_usbc_dsclen_3_14) 
);
defparam \u_usb_device_controller/usbc_dsclen_3_s8 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usbc_dsclen_4_s8  (
    .F(u_usb_device_controller_usbc_dsclen_4),
    .I0(u_usb_device_controller_usbc_dsclen_4_14),
    .I1(u_usb_device_controller_usbc_dsclen_4_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_4_s8 .INIT=16'h0305;
  LUT2 \u_usb_device_controller/usbc_dsclen_5_s8  (
    .F(u_usb_device_controller_usbc_dsclen_5),
    .I0(u_usb_device_controller_usbc_dsclen_0_28),
    .I1(u_usb_device_controller_usbc_dsclen_5_14) 
);
defparam \u_usb_device_controller/usbc_dsclen_5_s8 .INIT=4'h4;
  LUT2 \u_usb_device_controller/usbc_dsclen_7_s8  (
    .F(u_usb_device_controller_usbc_dsclen_7),
    .I0(u_usb_device_controller_usbc_dsclen_0_28),
    .I1(u_usb_device_controller_usbc_dsclen_7_14) 
);
defparam \u_usb_device_controller/usbc_dsclen_7_s8 .INIT=4'h4;
  LUT4 \u_usb_device_controller/descrom_start_0_s8  (
    .F(u_usb_device_controller_descrom_start_0),
    .I0(u_usb_device_controller_descrom_start_0_14),
    .I1(u_usb_device_controller_descrom_start_0_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_0_s8 .INIT=16'h030A;
  LUT4 \u_usb_device_controller/descrom_start_1_s8  (
    .F(u_usb_device_controller_descrom_start_1),
    .I0(u_usb_device_controller_descrom_start_1_14),
    .I1(u_usb_device_controller_descrom_start_1_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_1_s8 .INIT=16'h030A;
  LUT4 \u_usb_device_controller/descrom_start_2_s8  (
    .F(u_usb_device_controller_descrom_start_2),
    .I0(u_usb_device_controller_descrom_start_2_14),
    .I1(u_usb_device_controller_descrom_start_2_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_2_s8 .INIT=16'h030A;
  LUT4 \u_usb_device_controller/descrom_start_3_s8  (
    .F(u_usb_device_controller_descrom_start_3),
    .I0(u_usb_device_controller_descrom_start_3_14),
    .I1(u_usb_device_controller_descrom_start_3_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_3_s8 .INIT=16'h030A;
  LUT4 \u_usb_device_controller/descrom_start_4_s8  (
    .F(u_usb_device_controller_descrom_start_4),
    .I0(u_usb_device_controller_descrom_start_4_14),
    .I1(u_usb_device_controller_descrom_start_4_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_4_s8 .INIT=16'h030A;
  LUT4 \u_usb_device_controller/descrom_start_5_s8  (
    .F(u_usb_device_controller_descrom_start_5),
    .I0(u_usb_device_controller_descrom_start_5_14),
    .I1(u_usb_device_controller_descrom_start_5_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_5_s8 .INIT=16'h030A;
  LUT4 \u_usb_device_controller/descrom_start_6_s8  (
    .F(u_usb_device_controller_descrom_start_6),
    .I0(u_usb_device_controller_descrom_start_6_14),
    .I1(u_usb_device_controller_descrom_start_6_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_6_s8 .INIT=16'h030A;
  LUT4 \u_usb_device_controller/descrom_start_7_s8  (
    .F(u_usb_device_controller_descrom_start_7),
    .I0(u_usb_device_controller_descrom_start_7_14),
    .I1(u_usb_device_controller_descrom_start_7_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_7_s8 .INIT=16'h030A;
  LUT4 \u_usb_device_controller/descrom_start_8_s8  (
    .F(u_usb_device_controller_descrom_start_8),
    .I0(u_usb_device_controller_descrom_start_8_14),
    .I1(u_usb_device_controller_descrom_start_8_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_8_s8 .INIT=16'h030A;
  LUT4 \u_usb_device_controller/descrom_start_9_s8  (
    .F(u_usb_device_controller_descrom_start_9),
    .I0(u_usb_device_controller_descrom_start_9_14),
    .I1(u_usb_device_controller_descrom_start_9_15),
    .I2(u_usb_device_controller_usbc_dsclen_0_28),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/descrom_start_9_s8 .INIT=16'h030A;
  LUT2 \u_usb_device_controller/usb_transact_inst/txpop_o_d_s  (
    .F(u_usb_device_controller_usb_transact_inst_txpop_o_d),
    .I0(u_usb_device_controller_usb_transact_inst_txpop_o_d_9),
    .I1(u_usb_device_controller_usb_transact_inst_txpop_o_d_5) 
);
defparam \u_usb_device_controller/usb_transact_inst/txpop_o_d_s .INIT=4'h4;
  LUT3 \u_usb_device_controller/test_packet_inst/n315_s3  (
    .F(u_usb_device_controller_test_packet_inst_n315),
    .I0(u_usb_device_controller_test_packet_inst_n315_10),
    .I1(u_usb_device_controller_test_packet_inst_n312_9),
    .I2(u_usb_device_controller_test_packet_inst_n317_10) 
);
defparam \u_usb_device_controller/test_packet_inst/n315_s3 .INIT=8'hB0;
  LUT4 \u_usb_device_controller/test_packet_inst/n313_s3  (
    .F(u_usb_device_controller_test_packet_inst_n313),
    .I0(u_usb_device_controller_test_packet_inst_n133_6),
    .I1(u_usb_device_controller_test_packet_inst_test_data_val_9),
    .I2(u_usb_device_controller_test_packet_inst_n313_8),
    .I3(u_usb_device_controller_test_packet_inst_n317_10) 
);
defparam \u_usb_device_controller/test_packet_inst/n313_s3 .INIT=16'hF400;
  LUT3 \u_usb_device_controller/test_packet_inst/n316_s3  (
    .F(u_usb_device_controller_test_packet_inst_n316),
    .I0(u_usb_device_controller_test_packet_inst_n316_8),
    .I1(u_usb_device_controller_test_packet_inst_test_data_6),
    .I2(u_usb_device_controller_test_packet_inst_n312_10) 
);
defparam \u_usb_device_controller/test_packet_inst/n316_s3 .INIT=8'hE0;
  LUT4 \u_usb_device_controller/test_packet_inst/n314_s3  (
    .F(u_usb_device_controller_test_packet_inst_n314),
    .I0(u_usb_device_controller_test_packet_inst_n314_8),
    .I1(u_usb_device_controller_test_packet_inst_test_data_val_9),
    .I2(u_usb_device_controller_test_packet_inst_n313_8),
    .I3(u_usb_device_controller_test_packet_inst_n314_9) 
);
defparam \u_usb_device_controller/test_packet_inst/n314_s3 .INIT=16'hF400;
  LUT4 \u_usb_device_controller/u_usb_init/n211_s21  (
    .F(u_usb_device_controller_u_usb_init_n211),
    .I0(u_usb_device_controller_u_usb_init_s_state[3]),
    .I1(u_usb_device_controller_u_usb_init_s_state[2]),
    .I2(u_usb_device_controller_u_usb_init_s_state[1]),
    .I3(u_usb_device_controller_u_usb_init_s_state_0_4) 
);
defparam \u_usb_device_controller/u_usb_init/n211_s21 .INIT=16'h1FFF;
  LUT2 \u_usb_device_controller/usb_control_inst/n414_s1  (
    .F(u_usb_device_controller_usb_control_inst_n414),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n414_s1 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/n413_s1  (
    .F(u_usb_device_controller_usb_control_inst_n413),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n413_s1 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/n412_s1  (
    .F(u_usb_device_controller_usb_control_inst_n412),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n412_s1 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/n411_s1  (
    .F(u_usb_device_controller_usb_control_inst_n411),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n411_s1 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/n410_s1  (
    .F(u_usb_device_controller_usb_control_inst_n410),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n410_s1 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/n409_s1  (
    .F(u_usb_device_controller_usb_control_inst_n409),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n409_s1 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/n408_s1  (
    .F(u_usb_device_controller_usb_control_inst_n408),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n408_s1 .INIT=4'hE;
  LUT2 \u_usb_device_controller/usb_control_inst/n407_s1  (
    .F(u_usb_device_controller_usb_control_inst_n407),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n407_s1 .INIT=4'hE;
  LUT4 \u_usb_device_controller/u_usb_packet/n776_s1  (
    .F(u_usb_device_controller_u_usb_packet_n776),
    .I0(u_usb_device_controller_u_usb_packet_n776_6),
    .I1(u_usb_device_controller_u_usb_packet_n776_7),
    .I2(u_usb_device_controller_u_usb_packet_n776_8),
    .I3(u_usb_device_controller_u_usb_packet_n776_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n776_s1 .INIT=16'h96FF;
  LUT4 \u_usb_device_controller/u_usb_packet/n775_s1  (
    .F(u_usb_device_controller_u_usb_packet_n775),
    .I0(u_usb_device_controller_u_usb_packet_n775_6),
    .I1(u_usb_device_controller_u_usb_packet_n775_7),
    .I2(u_usb_device_controller_u_usb_packet_n775_8),
    .I3(u_usb_device_controller_u_usb_packet_n776_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n775_s1 .INIT=16'h69FF;
  LUT3 \u_usb_device_controller/u_usb_packet/n764_s1  (
    .F(u_usb_device_controller_u_usb_packet_n764),
    .I0(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I1(u_usb_device_controller_u_usb_packet_crc16_buf[4]),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n764_s1 .INIT=8'hFE;
  LUT4 \u_usb_device_controller/u_usb_packet/n761_s1  (
    .F(u_usb_device_controller_u_usb_packet_n761),
    .I0(u_usb_device_controller_u_usb_packet_n776_6),
    .I1(u_usb_device_controller_u_usb_packet_n776_8),
    .I2(u_usb_device_controller_u_usb_packet_n761_6),
    .I3(u_usb_device_controller_u_usb_packet_n776_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n761_s1 .INIT=16'h96FF;
  LUT4 \u_usb_device_controller/u_usb_init/n217_s27  (
    .F(u_usb_device_controller_u_usb_init_n217),
    .I0(u_usb_device_controller_u_usb_init_n217_37),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I2(u_usb_device_controller_u_usb_init_n217_38),
    .I3(u_usb_device_controller_u_usb_init_s_state[3]) 
);
defparam \u_usb_device_controller/u_usb_init/n217_s27 .INIT=16'hFF0B;
  LUT2 \u_usb_device_controller/utmi_opmode_o_d_1_s  (
    .F(u_usb_device_controller_utmi_opmode_o_d[1]),
    .I0(u_usb_device_controller_u_usb_init_usbi_opmode[1]),
    .I1(u_usb_device_controller_utmi_txvalid_o_d_8) 
);
defparam \u_usb_device_controller/utmi_opmode_o_d_1_s .INIT=4'hB;
  LUT2 \u_usb_device_controller/n1261_s1  (
    .F(u_usb_device_controller_n1261),
    .I0(txdat_len_i_d[10]),
    .I1(txdat_len_i_d[11]) 
);
defparam \u_usb_device_controller/n1261_s1 .INIT=4'hE;
  LUT4 \u_usb_device_controller/u_usb_packet/crc5_buf_4_s5  (
    .F(u_usb_device_controller_u_usb_packet_crc5_buf_4),
    .I0(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf_4_13),
    .I2(u_usb_device_controller_u_usb_packet_n784_18),
    .I3(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/u_usb_packet/crc5_buf_4_s5 .INIT=16'h00F8;
  LUT2 \u_usb_device_controller/usb_control_inst/s_answerptr_7_s6  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_7),
    .I0(u_usb_device_controller_usb_control_inst_s_answerptr_7_13),
    .I1(u_usb_device_controller_usb_control_inst_s_answerptr_7_8) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_7_s6 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s7  (
    .F(u_usb_device_controller_usb_control_inst_s_sendbyte_1),
    .I0(u_usb_device_controller_usb_control_inst_s_sendbyte_7_14),
    .I1(u_usb_device_controller_usb_control_inst_n2896_4),
    .I2(u_usb_device_controller_usb_control_inst_s_sendbyte_7_19),
    .I3(u_usb_device_controller_usb_control_inst_s_sendbyte_7_13) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s7 .INIT=16'h0B00;
  LUT3 \u_usb_device_controller/s_nyet_s4  (
    .F(u_usb_device_controller_s_nyet_9),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_n2393_9),
    .I2(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/s_nyet_s4 .INIT=8'hF8;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_sof_valid_s4  (
    .F(u_usb_device_controller_usb_transact_inst_s_sof_valid),
    .I0(u_usb_device_controller_usb_transact_inst_n1565_4),
    .I1(u_usb_device_controller_usb_transact_inst_n1041),
    .I2(u_usb_device_controller_usb_transact_inst_s_sof),
    .I3(u_usb_device_controller_usb_transact_inst_n1064_27) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sof_valid_s4 .INIT=16'hFF80;
  LUT2 \u_usb_device_controller/n1581_s1  (
    .F(u_usb_device_controller_n1581),
    .I0(u_usb_device_controller_s_endpt_rxrdy),
    .I1(u_usb_device_controller_rxact_o_d) 
);
defparam \u_usb_device_controller/n1581_s1 .INIT=4'h4;
  LUT2 \u_usb_device_controller/usb_control_inst/n1388_s4  (
    .F(u_usb_device_controller_usb_control_inst_n1388),
    .I0(inf_alter_i_d[1]),
    .I1(u_usb_device_controller_usb_control_inst_n1388_12) 
);
defparam \u_usb_device_controller/usb_control_inst/n1388_s4 .INIT=4'h8;
  LUT2 \u_usb_device_controller/usb_control_inst/n1387_s4  (
    .F(u_usb_device_controller_usb_control_inst_n1387),
    .I0(inf_alter_i_d[2]),
    .I1(u_usb_device_controller_usb_control_inst_n1388_12) 
);
defparam \u_usb_device_controller/usb_control_inst/n1387_s4 .INIT=4'h8;
  LUT2 \u_usb_device_controller/usb_control_inst/n1386_s4  (
    .F(u_usb_device_controller_usb_control_inst_n1386),
    .I0(inf_alter_i_d[3]),
    .I1(u_usb_device_controller_usb_control_inst_n1388_12) 
);
defparam \u_usb_device_controller/usb_control_inst/n1386_s4 .INIT=4'h8;
  LUT2 \u_usb_device_controller/usb_control_inst/n1385_s4  (
    .F(u_usb_device_controller_usb_control_inst_n1385),
    .I0(inf_alter_i_d[4]),
    .I1(u_usb_device_controller_usb_control_inst_n1388_12) 
);
defparam \u_usb_device_controller/usb_control_inst/n1385_s4 .INIT=4'h8;
  LUT2 \u_usb_device_controller/usb_control_inst/n1384_s4  (
    .F(u_usb_device_controller_usb_control_inst_n1384),
    .I0(inf_alter_i_d[5]),
    .I1(u_usb_device_controller_usb_control_inst_n1388_12) 
);
defparam \u_usb_device_controller/usb_control_inst/n1384_s4 .INIT=4'h8;
  LUT2 \u_usb_device_controller/usb_control_inst/n1383_s4  (
    .F(u_usb_device_controller_usb_control_inst_n1383),
    .I0(inf_alter_i_d[6]),
    .I1(u_usb_device_controller_usb_control_inst_n1388_12) 
);
defparam \u_usb_device_controller/usb_control_inst/n1383_s4 .INIT=4'h8;
  LUT2 \u_usb_device_controller/usb_control_inst/n1382_s4  (
    .F(u_usb_device_controller_usb_control_inst_n1382),
    .I0(inf_alter_i_d[7]),
    .I1(u_usb_device_controller_usb_control_inst_n1388_12) 
);
defparam \u_usb_device_controller/usb_control_inst/n1382_s4 .INIT=4'h8;
  LUT3 \u_usb_device_controller/usb_control_inst/n1617_s1  (
    .F(u_usb_device_controller_usb_control_inst_n1617),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[6]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[7]),
    .I2(u_usb_device_controller_usb_control_inst_n1670_39) 
);
defparam \u_usb_device_controller/usb_control_inst/n1617_s1 .INIT=8'h60;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1136_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1136),
    .I0(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[9]),
    .I2(u_usb_device_controller_usb_transact_inst_n1138_39) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1136_s19 .INIT=8'h14;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1133_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1133),
    .I0(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[10]),
    .I2(u_usb_device_controller_usb_transact_inst_n1133_26) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1133_s19 .INIT=8'h14;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1130_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1130),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[10]),
    .I1(u_usb_device_controller_usb_transact_inst_n1133_26),
    .I2(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[11]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1130_s19 .INIT=16'h0B04;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1127_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1127),
    .I0(u_usb_device_controller_usb_transact_inst_n1133_26),
    .I1(u_usb_device_controller_usb_transact_inst_n1127_26),
    .I2(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[12]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1127_s19 .INIT=16'h0708;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1124_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1124),
    .I0(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[13]),
    .I2(u_usb_device_controller_usb_transact_inst_n1124_28) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1124_s19 .INIT=8'h14;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1121_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1121),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[13]),
    .I1(u_usb_device_controller_usb_transact_inst_n1124_28),
    .I2(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[14]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1121_s19 .INIT=16'h0B04;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1118_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1118),
    .I0(u_usb_device_controller_usb_transact_inst_n1124_28),
    .I1(u_usb_device_controller_usb_transact_inst_n1118_26),
    .I2(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[15]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1118_s19 .INIT=16'h0708;
  LUT4 \u_usb_device_controller/n1609_s14  (
    .F(u_usb_device_controller_n1609),
    .I0(u_usb_device_controller_s_bufptr[2]),
    .I1(u_usb_device_controller_n1611_21),
    .I2(u_usb_device_controller_n1613_21),
    .I3(u_usb_device_controller_s_bufptr[3]) 
);
defparam \u_usb_device_controller/n1609_s14 .INIT=16'h0708;
  LUT4 \u_usb_device_controller/n1605_s14  (
    .F(u_usb_device_controller_n1605),
    .I0(u_usb_device_controller_s_bufptr[4]),
    .I1(u_usb_device_controller_n1607_23),
    .I2(u_usb_device_controller_n1613_21),
    .I3(u_usb_device_controller_s_bufptr[5]) 
);
defparam \u_usb_device_controller/n1605_s14 .INIT=16'h0708;
  LUT4 \u_usb_device_controller/n1603_s14  (
    .F(u_usb_device_controller_n1603),
    .I0(u_usb_device_controller_n1607_23),
    .I1(u_usb_device_controller_n1603_21),
    .I2(u_usb_device_controller_n1613_21),
    .I3(u_usb_device_controller_s_bufptr[6]) 
);
defparam \u_usb_device_controller/n1603_s14 .INIT=16'h0708;
  LUT4 \u_usb_device_controller/n1599_s14  (
    .F(u_usb_device_controller_n1599),
    .I0(u_usb_device_controller_s_bufptr[7]),
    .I1(u_usb_device_controller_n1601_23),
    .I2(u_usb_device_controller_n1613_21),
    .I3(u_usb_device_controller_s_bufptr[8]) 
);
defparam \u_usb_device_controller/n1599_s14 .INIT=16'h0708;
  LUT4 \u_usb_device_controller/n1597_s14  (
    .F(u_usb_device_controller_n1597),
    .I0(u_usb_device_controller_n1601_23),
    .I1(u_usb_device_controller_n1597_21),
    .I2(u_usb_device_controller_n1613_21),
    .I3(u_usb_device_controller_s_bufptr[9]) 
);
defparam \u_usb_device_controller/n1597_s14 .INIT=16'h0708;
  LUT4 \u_usb_device_controller/n1593_s15  (
    .F(u_usb_device_controller_n1593),
    .I0(u_usb_device_controller_s_bufptr[10]),
    .I1(u_usb_device_controller_n1595_23),
    .I2(u_usb_device_controller_n1613_21),
    .I3(u_usb_device_controller_s_bufptr[11]) 
);
defparam \u_usb_device_controller/n1593_s15 .INIT=16'h0708;
  LUT3 \u_usb_device_controller/u_usb_packet/n579_s12  (
    .F(u_usb_device_controller_u_usb_packet_n579),
    .I0(u_usb_device_controller_u_usb_packet_n579_19),
    .I1(u_usb_device_controller_u_usb_packet_n579_20),
    .I2(u_usb_device_controller_u_usb_packet_n784_18) 
);
defparam \u_usb_device_controller/u_usb_packet/n579_s12 .INIT=8'hF8;
  LUT4 \u_usb_device_controller/u_usb_packet/n577_s12  (
    .F(u_usb_device_controller_u_usb_packet_n577),
    .I0(u_usb_device_controller_u_usb_packet_n784_18),
    .I1(u_usb_device_controller_u_usb_packet_n577_19),
    .I2(u_usb_device_controller_u_usb_packet_n577_20),
    .I3(u_usb_device_controller_u_usb_packet_n579_20) 
);
defparam \u_usb_device_controller/u_usb_packet/n577_s12 .INIT=16'hBEAA;
  LUT4 \u_usb_device_controller/u_usb_packet/n575_s12  (
    .F(u_usb_device_controller_u_usb_packet_n575),
    .I0(u_usb_device_controller_u_usb_packet_n784_18),
    .I1(u_usb_device_controller_u_usb_packet_n575_19),
    .I2(u_usb_device_controller_u_usb_packet_n577_20),
    .I3(u_usb_device_controller_u_usb_packet_n579_20) 
);
defparam \u_usb_device_controller/u_usb_packet/n575_s12 .INIT=16'hBEAA;
  LUT4 \u_usb_device_controller/u_usb_packet/n573_s12  (
    .F(u_usb_device_controller_u_usb_packet_n573),
    .I0(u_usb_device_controller_u_usb_packet_n784_18),
    .I1(u_usb_device_controller_u_usb_packet_n573_19),
    .I2(u_usb_device_controller_u_usb_packet_n577_19),
    .I3(u_usb_device_controller_u_usb_packet_n579_20) 
);
defparam \u_usb_device_controller/u_usb_packet/n573_s12 .INIT=16'hBEAA;
  LUT3 \u_usb_device_controller/u_usb_packet/n571_s12  (
    .F(u_usb_device_controller_u_usb_packet_n571),
    .I0(u_usb_device_controller_u_usb_packet_n571_19),
    .I1(u_usb_device_controller_u_usb_packet_n579_20),
    .I2(u_usb_device_controller_u_usb_packet_n784_18) 
);
defparam \u_usb_device_controller/u_usb_packet/n571_s12 .INIT=8'hF8;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_7_s1  (
    .F(u_usb_device_controller_utmi_dataout_o_d_7),
    .I0(u_usb_device_controller_test_packet_inst_test_data_Z[7]),
    .I1(u_usb_device_controller_u_usb_packet_usbp_dataout_o[7]),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_7),
    .I3(u_usb_device_controller_utmi_txvalid_o_d_6) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_7_s1 .INIT=16'h0A0C;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_6_s0  (
    .F(u_usb_device_controller_utmi_dataout_o_d_6),
    .I0(u_usb_device_controller_test_packet_inst_test_data_Z[6]),
    .I1(u_usb_device_controller_u_usb_packet_usbp_dataout_o[6]),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_7),
    .I3(u_usb_device_controller_utmi_txvalid_o_d_6) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_6_s0 .INIT=16'h0A0C;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_5_s0  (
    .F(u_usb_device_controller_utmi_dataout_o_d_5),
    .I0(u_usb_device_controller_test_packet_inst_test_data_Z[5]),
    .I1(u_usb_device_controller_u_usb_packet_usbp_dataout_o[5]),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_7),
    .I3(u_usb_device_controller_utmi_txvalid_o_d_6) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_5_s0 .INIT=16'h0A0C;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_4_s0  (
    .F(u_usb_device_controller_utmi_dataout_o_d_4),
    .I0(u_usb_device_controller_test_packet_inst_test_data_Z[4]),
    .I1(u_usb_device_controller_u_usb_packet_usbp_dataout_o[4]),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_7),
    .I3(u_usb_device_controller_utmi_txvalid_o_d_6) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_4_s0 .INIT=16'h0A0C;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_3_s0  (
    .F(u_usb_device_controller_utmi_dataout_o_d_3),
    .I0(u_usb_device_controller_test_packet_inst_test_data_Z[3]),
    .I1(u_usb_device_controller_u_usb_packet_usbp_dataout_o[3]),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_7),
    .I3(u_usb_device_controller_utmi_txvalid_o_d_6) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_3_s0 .INIT=16'h0A0C;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_2_s0  (
    .F(u_usb_device_controller_utmi_dataout_o_d_2),
    .I0(u_usb_device_controller_test_packet_inst_test_data_Z[2]),
    .I1(u_usb_device_controller_u_usb_packet_usbp_dataout_o[2]),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_7),
    .I3(u_usb_device_controller_utmi_txvalid_o_d_6) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_2_s0 .INIT=16'h0A0C;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_1_s0  (
    .F(u_usb_device_controller_utmi_dataout_o_d_1),
    .I0(u_usb_device_controller_test_packet_inst_test_data_Z[1]),
    .I1(u_usb_device_controller_u_usb_packet_usbp_dataout_o[1]),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_7),
    .I3(u_usb_device_controller_utmi_txvalid_o_d_6) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_1_s0 .INIT=16'h0A0C;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_0_s0  (
    .F(u_usb_device_controller_utmi_dataout_o_d_0),
    .I0(u_usb_device_controller_utmi_dataout_o_d_7_10),
    .I1(u_usb_device_controller_utmi_dataout_o_d_0_4),
    .I2(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I3(u_usb_device_controller_utmi_dataout_o_d_0_5) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_0_s0 .INIT=16'hF3A0;
  LUT2 \u_usb_device_controller/rxact_o_d_s0  (
    .F(u_usb_device_controller_rxact_o_d_3),
    .I0(u_usb_device_controller_cur_state[3]),
    .I1(u_usb_device_controller_cur_state[2]) 
);
defparam \u_usb_device_controller/rxact_o_d_s0 .INIT=4'h4;
  LUT4 \u_usb_device_controller/n2339_s1  (
    .F(u_usb_device_controller_n2339_4),
    .I0(txdat_len_i_d[0]),
    .I1(txdat_len_i_d[1]),
    .I2(u_usb_device_controller_n2339_5),
    .I3(u_usb_device_controller_n2339_6) 
);
defparam \u_usb_device_controller/n2339_s1 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/n1585_s1  (
    .F(u_usb_device_controller_n1585_4),
    .I0(u_usb_device_controller_cur_state[2]),
    .I1(u_usb_device_controller_cur_state[3]) 
);
defparam \u_usb_device_controller/n1585_s1 .INIT=4'h1;
  LUT2 \u_usb_device_controller/setup_o_d_s0  (
    .F(u_usb_device_controller_setup_o_d_3),
    .I0(u_usb_device_controller_cur_state[0]),
    .I1(u_usb_device_controller_cur_state[1]) 
);
defparam \u_usb_device_controller/setup_o_d_s0 .INIT=4'h1;
  LUT4 \u_usb_device_controller/n2024_s1  (
    .F(u_usb_device_controller_n2024_4),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[6]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I2(u_usb_device_controller_n2024_5),
    .I3(u_usb_device_controller_n2024_6) 
);
defparam \u_usb_device_controller/n2024_s1 .INIT=16'h4000;
  LUT3 \u_usb_device_controller/test_packet_inst/n127_s3  (
    .F(u_usb_device_controller_test_packet_inst_n127_6),
    .I0(u_usb_device_controller_test_packet_inst_cnt[8]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[9]),
    .I2(u_usb_device_controller_test_packet_inst_n129_6) 
);
defparam \u_usb_device_controller/test_packet_inst/n127_s3 .INIT=8'h80;
  LUT3 \u_usb_device_controller/test_packet_inst/n127_s4  (
    .F(u_usb_device_controller_test_packet_inst_n127_7),
    .I0(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I1(u_usb_device_controller_test_packet_inst_n378_4),
    .I2(u_usb_device_controller_test_packet_inst_test_en_dect) 
);
defparam \u_usb_device_controller/test_packet_inst/n127_s4 .INIT=8'h10;
  LUT3 \u_usb_device_controller/test_packet_inst/n129_s3  (
    .F(u_usb_device_controller_test_packet_inst_n129_6),
    .I0(u_usb_device_controller_test_packet_inst_cnt[6]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[7]),
    .I2(u_usb_device_controller_test_packet_inst_n131_8) 
);
defparam \u_usb_device_controller/test_packet_inst/n129_s3 .INIT=8'h80;
  LUT4 \u_usb_device_controller/test_packet_inst/n130_s3  (
    .F(u_usb_device_controller_test_packet_inst_n130_6),
    .I0(u_usb_device_controller_test_packet_inst_cnt[7]),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_test_packet_inst_n130_7),
    .I3(u_usb_device_controller_test_packet_inst_n127_7) 
);
defparam \u_usb_device_controller/test_packet_inst/n130_s3 .INIT=16'h00BF;
  LUT3 \u_usb_device_controller/test_packet_inst/n133_s3  (
    .F(u_usb_device_controller_test_packet_inst_n133_6),
    .I0(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[2]) 
);
defparam \u_usb_device_controller/test_packet_inst/n133_s3 .INIT=8'h80;
  LUT2 \u_usb_device_controller/test_packet_inst/n133_s4  (
    .F(u_usb_device_controller_test_packet_inst_n133_7),
    .I0(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[4]) 
);
defparam \u_usb_device_controller/test_packet_inst/n133_s4 .INIT=4'h8;
  LUT4 \u_usb_device_controller/test_packet_inst/n378_s1  (
    .F(u_usb_device_controller_test_packet_inst_n378_4),
    .I0(u_usb_device_controller_test_packet_inst_n378_5),
    .I1(u_usb_device_controller_test_packet_inst_n378_8),
    .I2(u_usb_device_controller_test_packet_inst_cnt[10]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[11]) 
);
defparam \u_usb_device_controller/test_packet_inst/n378_s1 .INIT=16'hD000;
  LUT2 \u_usb_device_controller/u_usb_init/n414_s1  (
    .F(u_usb_device_controller_u_usb_init_n414_4),
    .I0(u_usb_device_controller_u_usb_init_s_state[2]),
    .I1(u_usb_device_controller_u_usb_init_s_state[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n414_s1 .INIT=4'h4;
  LUT2 \u_usb_device_controller/u_usb_packet/n782_s1  (
    .F(u_usb_device_controller_u_usb_packet_n782_4),
    .I0(u_usb_device_controller_u_usb_packet_n782_6),
    .I1(u_usb_device_controller_u_usb_packet_n782_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n782_s1 .INIT=4'h4;
  LUT2 \u_usb_device_controller/u_usb_packet/n782_s2  (
    .F(u_usb_device_controller_u_usb_packet_n782_5),
    .I0(u_usb_device_controller_u_usb_packet_n782_8),
    .I1(u_usb_device_controller_u_usb_packet_n782_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n782_s2 .INIT=4'h1;
  LUT4 \u_usb_device_controller/u_usb_packet/n784_s1  (
    .F(u_usb_device_controller_u_usb_packet_n784_4),
    .I0(u_usb_device_controller_u_usb_packet_n622),
    .I1(u_usb_device_controller_u_usb_packet_crc16_buf[14]),
    .I2(u_usb_device_controller_u_usb_packet_n784_7),
    .I3(u_usb_device_controller_u_usb_packet_n784_8) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s1 .INIT=16'h0D00;
  LUT3 \u_usb_device_controller/u_usb_packet/n784_s3  (
    .F(u_usb_device_controller_u_usb_packet_n784_6),
    .I0(u_usb_device_controller_u_usb_packet_n328_10),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[1]),
    .I2(u_usb_device_controller_u_usb_packet_n784_16) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s3 .INIT=8'hAC;
  LUT3 \u_usb_device_controller/u_usb_packet/n785_s1  (
    .F(u_usb_device_controller_u_usb_packet_n785_4),
    .I0(u_usb_device_controller_u_usb_packet_n785_6),
    .I1(u_usb_device_controller_u_usb_packet_n328_11),
    .I2(u_usb_device_controller_u_usb_packet_n785_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n785_s1 .INIT=8'h70;
  LUT3 \u_usb_device_controller/u_usb_packet/n785_s2  (
    .F(u_usb_device_controller_u_usb_packet_n785_5),
    .I0(u_usb_device_controller_u_usb_packet_n328_11),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[0]),
    .I2(u_usb_device_controller_u_usb_packet_n784_16) 
);
defparam \u_usb_device_controller/u_usb_packet/n785_s2 .INIT=8'hAC;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s1  (
    .F(u_usb_device_controller_u_usb_packet_n912_4),
    .I0(u_usb_device_controller_u_usb_packet_n774_6),
    .I1(u_usb_device_controller_u_usb_packet_n764),
    .I2(u_usb_device_controller_u_usb_packet_n770_6),
    .I3(u_usb_device_controller_u_usb_packet_n912_8) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s1 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s2  (
    .F(u_usb_device_controller_u_usb_packet_n912_5),
    .I0(u_usb_device_controller_u_usb_packet_n912_9),
    .I1(u_usb_device_controller_u_usb_packet_n767_6),
    .I2(u_usb_device_controller_u_usb_packet_n912_10),
    .I3(u_usb_device_controller_u_usb_packet_n771_6) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s2 .INIT=16'h0001;
  LUT2 \u_usb_device_controller/u_usb_packet/n912_s3  (
    .F(u_usb_device_controller_u_usb_packet_n912_6),
    .I0(u_usb_device_controller_u_usb_packet_n774_7),
    .I1(u_usb_device_controller_u_usb_packet_n771_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s3 .INIT=4'h1;
  LUT3 \u_usb_device_controller/u_usb_packet/n912_s4  (
    .F(u_usb_device_controller_u_usb_packet_n912_7),
    .I0(u_usb_device_controller_u_usb_packet_n912_11),
    .I1(u_usb_device_controller_u_usb_packet_n912_12),
    .I2(u_usb_device_controller_u_usb_packet_n912_13) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s4 .INIT=8'hD0;
  LUT4 \u_usb_device_controller/u_usb_packet/n920_s1  (
    .F(u_usb_device_controller_u_usb_packet_n920_4),
    .I0(u_usb_device_controller_u_usb_packet_n920_6),
    .I1(u_usb_device_controller_u_usb_packet_s_txready),
    .I2(u_usb_device_controller_u_usb_packet_n626),
    .I3(u_usb_device_controller_u_usb_packet_n920_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n920_s1 .INIT=16'h0D00;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1041_s1  (
    .F(u_usb_device_controller_usb_transact_inst_n1041_4),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[5]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[6]),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[7]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1041_s1 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1041_s3  (
    .F(u_usb_device_controller_usb_transact_inst_n1041_6),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[0]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[1]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[3]),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[2]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1041_s3 .INIT=16'h0100;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1565_s1  (
    .F(u_usb_device_controller_usb_transact_inst_n1565_4),
    .I0(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I1(u_usb_device_controller_u_usb_packet_s_rxvalid) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1565_s1 .INIT=4'h8;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1565_s2  (
    .F(u_usb_device_controller_usb_transact_inst_n1565_5),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1565_s2 .INIT=4'h8;
  LUT4 \u_usb_device_controller/usb_control_inst/n1629_s1  (
    .F(u_usb_device_controller_usb_control_inst_n1629_4),
    .I0(u_usb_device_controller_usb_control_inst_s_state[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[1]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[2]),
    .I3(u_usb_device_controller_usb_control_inst_s_state[3]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1629_s1 .INIT=16'h0001;
  LUT3 \u_usb_device_controller/usb_control_inst/n1629_s2  (
    .F(u_usb_device_controller_usb_control_inst_n1629_5),
    .I0(u_usb_device_controller_usb_control_inst_s_state[7]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[8]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[9]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1629_s2 .INIT=8'h01;
  LUT3 \u_usb_device_controller/usb_control_inst/n1629_s3  (
    .F(u_usb_device_controller_usb_control_inst_n1629_6),
    .I0(u_usb_device_controller_usb_control_inst_s_state[5]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[4]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1629_s3 .INIT=8'h10;
  LUT2 \u_usb_device_controller/usb_control_inst/n2896_s1  (
    .F(u_usb_device_controller_usb_control_inst_n2896_4),
    .I0(u_usb_device_controller_usb_transact_inst_s_setup_2),
    .I1(u_usb_device_controller_usb_control_inst_n2896_9) 
);
defparam \u_usb_device_controller/usb_control_inst/n2896_s1 .INIT=4'h4;
  LUT2 \u_usb_device_controller/usb_control_inst/n2896_s2  (
    .F(u_usb_device_controller_usb_control_inst_n2896_5),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n2896_s2 .INIT=4'h4;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s20  (
    .F(u_usb_device_controller_u_usb_init_n212_28),
    .I0(u_usb_device_controller_u_usb_init_n212_57),
    .I1(u_usb_device_controller_u_usb_init_s_opmode_1),
    .I2(u_usb_device_controller_u_usb_init_n212_33),
    .I3(u_usb_device_controller_u_usb_init_n212_65) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s20 .INIT=16'h0BBB;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s21  (
    .F(u_usb_device_controller_u_usb_init_n212_29),
    .I0(u_usb_device_controller_u_usb_init_n212_35),
    .I1(u_usb_device_controller_u_usb_init_n212_59),
    .I2(u_usb_device_controller_u_usb_init_n212_37),
    .I3(u_usb_device_controller_u_usb_init_s_state[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s21 .INIT=16'hBB0F;
  LUT2 \u_usb_device_controller/u_usb_init/n212_s23  (
    .F(u_usb_device_controller_u_usb_init_n212_31),
    .I0(u_usb_device_controller_u_usb_init_s_state[3]),
    .I1(u_usb_device_controller_u_usb_init_s_state[2]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s23 .INIT=4'h4;
  LUT4 \u_usb_device_controller/u_usb_init/n215_s45  (
    .F(u_usb_device_controller_u_usb_init_n215_52),
    .I0(u_usb_device_controller_u_usb_init_n215_65),
    .I1(u_usb_device_controller_u_usb_init_n218),
    .I2(u_usb_device_controller_u_usb_init_n215_69),
    .I3(u_usb_device_controller_u_usb_init_n215_57) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s45 .INIT=16'h0B00;
  LUT4 \u_usb_device_controller/u_usb_init/n216_s43  (
    .F(u_usb_device_controller_u_usb_init_n216_49),
    .I0(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .I1(u_usb_device_controller_u_usb_init_s_linestate[1]),
    .I2(u_usb_device_controller_u_usb_init_n216_52),
    .I3(u_usb_device_controller_u_usb_init_n216_53) 
);
defparam \u_usb_device_controller/u_usb_init/n216_s43 .INIT=16'h004F;
  LUT4 \u_usb_device_controller/u_usb_init/n216_s45  (
    .F(u_usb_device_controller_u_usb_init_n216_51),
    .I0(u_usb_device_controller_u_usb_init_n215_53),
    .I1(u_usb_device_controller_u_usb_init_n215_54),
    .I2(u_usb_device_controller_u_usb_init_s_state[1]),
    .I3(u_usb_device_controller_u_usb_init_s_state[3]) 
);
defparam \u_usb_device_controller/u_usb_init/n216_s45 .INIT=16'hF400;
  LUT4 \u_usb_device_controller/usb_control_inst/n435_s12  (
    .F(u_usb_device_controller_usb_control_inst_n435_16),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I1(u_usb_device_controller_usb_control_inst_n435_18),
    .I2(u_usb_device_controller_usb_control_inst_n435_19),
    .I3(u_usb_device_controller_usb_control_inst_s_setupptr[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n435_s12 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/usb_control_inst/n435_s13  (
    .F(u_usb_device_controller_usb_control_inst_n435_17),
    .I0(u_usb_device_controller_usb_control_inst_n435_20),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I3(u_usb_device_controller_usb_control_inst_s_setupptr[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n435_s13 .INIT=16'h0D00;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s6  (
    .F(u_usb_device_controller_u_usb_packet_n328_10),
    .I0(u_usb_device_controller_u_usb_packet_n328_12),
    .I1(u_usb_device_controller_u_usb_packet_n328_13),
    .I2(u_usb_device_controller_u_usb_packet_n328_14),
    .I3(u_usb_device_controller_u_usb_packet_n328_31) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s6 .INIT=16'h004F;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s7  (
    .F(u_usb_device_controller_u_usb_packet_n328_11),
    .I0(u_usb_device_controller_u_usb_packet_n328_16),
    .I1(u_usb_device_controller_u_usb_packet_n328_17),
    .I2(u_usb_device_controller_u_usb_packet_n328_27),
    .I3(u_usb_device_controller_u_usb_packet_n328_29) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s7 .INIT=16'h008F;
  LUT4 \u_usb_device_controller/usb_control_inst/n1836_s5  (
    .F(u_usb_device_controller_usb_control_inst_n1836_8),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .I2(u_usb_device_controller_usb_control_inst_n1836_10),
    .I3(u_usb_device_controller_usb_control_inst_n2902_5) 
);
defparam \u_usb_device_controller/usb_control_inst/n1836_s5 .INIT=16'h0100;
  LUT3 \u_usb_device_controller/usb_control_inst/n1837_s3  (
    .F(u_usb_device_controller_usb_control_inst_n1837_6),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1837_s3 .INIT=8'h40;
  LUT3 \u_usb_device_controller/usb_control_inst/n1837_s4  (
    .F(u_usb_device_controller_usb_control_inst_n1837_7),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1837_s4 .INIT=8'h10;
  LUT2 \u_usb_device_controller/usb_control_inst/n2067_s3  (
    .F(u_usb_device_controller_usb_control_inst_n2067_6),
    .I0(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I1(u_usb_device_controller_usb_control_inst_n1836_15) 
);
defparam \u_usb_device_controller/usb_control_inst/n2067_s3 .INIT=4'h4;
  LUT2 \u_usb_device_controller/usb_control_inst/n2067_s4  (
    .F(u_usb_device_controller_usb_control_inst_n2067_7),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n2067_s4 .INIT=4'h8;
  LUT4 \u_usb_device_controller/u_usb_packet/n800_s3  (
    .F(u_usb_device_controller_u_usb_packet_n800_6),
    .I0(u_usb_device_controller_u_usb_packet_s_state[4]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[6]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[5]),
    .I3(u_usb_device_controller_u_usb_packet_n800_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n800_s3 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/rxdat_d0_7_s4  (
    .F(u_usb_device_controller_rxdat_d0_7_9),
    .I0(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I1(u_usb_device_controller_usb_transact_inst_s_out_valid) 
);
defparam \u_usb_device_controller/rxdat_d0_7_s4 .INIT=4'h4;
  LUT3 \u_usb_device_controller/rxdat_d0_7_s5  (
    .F(u_usb_device_controller_rxdat_d0_7_10),
    .I0(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I1(u_usb_device_controller_usb_transact_inst_s_setup_2),
    .I2(u_usb_device_controller_setup_o_d) 
);
defparam \u_usb_device_controller/rxdat_d0_7_s5 .INIT=8'hB0;
  LUT2 \u_usb_device_controller/u_usb_init/s_opmode_1_s4  (
    .F(u_usb_device_controller_u_usb_init_s_opmode_1),
    .I0(u_usb_device_controller_u_usb_init_s_state[1]),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4) 
);
defparam \u_usb_device_controller/u_usb_init/s_opmode_1_s4 .INIT=4'h1;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_3_s4  (
    .F(u_usb_device_controller_u_usb_init_s_state_3),
    .I0(u_usb_device_controller_u_usb_init_n212_39),
    .I1(u_usb_device_controller_u_usb_init_n414_4),
    .I2(u_usb_device_controller_u_usb_init_s_state_3_11),
    .I3(u_usb_device_controller_u_usb_init_s_state_2_14) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s4 .INIT=16'h7F00;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_3_s5  (
    .F(u_usb_device_controller_u_usb_init_s_state_3_10),
    .I0(u_usb_device_controller_u_usb_init_n214),
    .I1(u_usb_device_controller_u_usb_init_s_state_3_12),
    .I2(u_usb_device_controller_u_usb_init_n212_63),
    .I3(u_usb_device_controller_u_usb_init_s_state_2_18) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s5 .INIT=16'h000D;
  LUT4 \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s4  (
    .F(u_usb_device_controller_u_usb_init_s_chirpcnt_2_8),
    .I0(u_usb_device_controller_u_usb_init_s_chirpcnt_2_9),
    .I1(u_usb_device_controller_u_usb_init_n212_59),
    .I2(u_usb_device_controller_u_usb_init_s_chirpcnt_2_10),
    .I3(u_usb_device_controller_u_usb_init_s_state[1]) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s4 .INIT=16'h770F;
  LUT3 \u_usb_device_controller/usb_control_inst/s_answerlen_7_s3  (
    .F(u_usb_device_controller_usb_control_inst_s_answerlen_7_7),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen_7_11),
    .I2(u_usb_device_controller_usb_control_inst_s_answerlen_7_13) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerlen_7_s3 .INIT=8'h80;
  LUT4 \u_usb_device_controller/u_usb_packet/n615_s38  (
    .F(u_usb_device_controller_u_usb_packet_n615_42),
    .I0(u_usb_device_controller_u_usb_packet_n800_6),
    .I1(u_usb_device_controller_u_usb_packet_n615_44),
    .I2(u_usb_device_controller_u_usb_packet_n615_45),
    .I3(u_usb_device_controller_u_usb_packet_n615_46) 
);
defparam \u_usb_device_controller/u_usb_packet/n615_s38 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/u_usb_packet/s_dataout_7_s5  (
    .F(u_usb_device_controller_u_usb_packet_s_dataout_7_9),
    .I0(u_usb_device_controller_u_usb_packet_s_state[0]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[1]),
    .I2(u_usb_device_controller_u_usb_packet_n784_9),
    .I3(u_usb_device_controller_u_usb_packet_n784_10) 
);
defparam \u_usb_device_controller/u_usb_packet/s_dataout_7_s5 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1080_s41  (
    .F(u_usb_device_controller_usb_transact_inst_n1080),
    .I0(u_usb_device_controller_usb_transact_inst_n1041_4),
    .I1(u_usb_device_controller_usb_transact_inst_n1041_8),
    .I2(u_usb_device_controller_usb_transact_inst_n1080_48) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1080_s41 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1080_s42  (
    .F(u_usb_device_controller_usb_transact_inst_n1080_46),
    .I0(u_usb_device_controller_usb_transact_inst_n1080_49),
    .I1(u_usb_device_controller_usb_transact_inst_n1080_53),
    .I2(u_usb_device_controller_usb_transact_inst_n1095_45),
    .I3(u_usb_device_controller_usb_transact_inst_n1072_18) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1080_s42 .INIT=16'h000B;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1064_s11  (
    .F(u_usb_device_controller_usb_transact_inst_n1064_16),
    .I0(u_usb_device_controller_usb_transact_inst_n1157_26),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_27),
    .I2(u_usb_device_controller_usb_transact_inst_n1041_4),
    .I3(u_usb_device_controller_usb_transact_inst_n1064_20) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1064_s11 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1074_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1074_22),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[0]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[1]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[3]),
    .I3(u_usb_device_controller_usb_transact_inst_n1074_25) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1074_s17 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1072_s12  (
    .F(u_usb_device_controller_usb_transact_inst_n1072_18),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[7]),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_27),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_28),
    .I3(u_usb_device_controller_usb_transact_inst_n1072_21) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1072_s12 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1072_s13  (
    .F(u_usb_device_controller_usb_transact_inst_n1072_19),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[11]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[12]),
    .I3(u_usb_device_controller_usb_transact_inst_n1080_53) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1072_s13 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1138_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_24),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[12]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[11]),
    .I3(u_usb_device_controller_usb_transact_inst_n1080_53) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s19 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1138_s20  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_25),
    .I0(u_usb_device_controller_usb_transact_inst_txpop_o_d_5),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I2(u_usb_device_controller_usb_transact_inst_n1064_16) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s20 .INIT=8'h01;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1157_s20  (
    .F(u_usb_device_controller_usb_transact_inst_n1157_26),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[9]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1157_s20 .INIT=4'h1;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1157_s21  (
    .F(u_usb_device_controller_usb_transact_inst_n1157_27),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[0]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[1]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[2]),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[3]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1157_s21 .INIT=16'h0001;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1157_s22  (
    .F(u_usb_device_controller_usb_transact_inst_n1157_28),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[10]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[11]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[12]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1157_s22 .INIT=8'h01;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1157_s23  (
    .F(u_usb_device_controller_usb_transact_inst_n1157_29),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[5]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[6]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[7]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1157_s23 .INIT=16'h0110;
  LUT3 \u_usb_device_controller/usb_control_inst/n1670_s35  (
    .F(u_usb_device_controller_usb_control_inst_n1670_39),
    .I0(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_11) 
);
defparam \u_usb_device_controller/usb_control_inst/n1670_s35 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1670_s36  (
    .F(u_usb_device_controller_usb_control_inst_n1670_40),
    .I0(u_usb_device_controller_usb_control_inst_n1629),
    .I1(u_usb_device_controller_usb_control_inst_n1678_40),
    .I2(u_usb_device_controller_usb_control_inst_n1686_39),
    .I3(u_usb_device_controller_usb_control_inst_n1684_39) 
);
defparam \u_usb_device_controller/usb_control_inst/n1670_s36 .INIT=16'h0001;
  LUT3 \u_usb_device_controller/usb_control_inst/n1670_s37  (
    .F(u_usb_device_controller_usb_control_inst_n1670_41),
    .I0(u_usb_device_controller_usb_control_inst_s_answerptr_5_10),
    .I1(u_usb_device_controller_usb_control_inst_n1670_43),
    .I2(u_usb_device_controller_usb_control_inst_s_interface_set_8) 
);
defparam \u_usb_device_controller/usb_control_inst/n1670_s37 .INIT=8'h01;
  LUT3 \u_usb_device_controller/usb_control_inst/s_answerptr_7_s7  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_7_11),
    .I0(u_usb_device_controller_usb_control_inst_s_state[7]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[8]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_14) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_7_s7 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_control_inst/s_answerptr_7_s8  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_7_12),
    .I0(u_usb_device_controller_usb_control_inst_s_state[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[1]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_15) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_7_s8 .INIT=8'h40;
  LUT3 \u_usb_device_controller/usb_control_inst/s_answerptr_5_s7  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_5_10),
    .I0(u_usb_device_controller_usb_control_inst_n1629_4),
    .I1(u_usb_device_controller_usb_control_inst_n1629_5),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_5_12) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_5_s7 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s9  (
    .F(u_usb_device_controller_usb_control_inst_s_sendbyte_7_13),
    .I0(u_usb_device_controller_usb_control_inst_n2896_4),
    .I1(u_usb_device_controller_usb_control_inst_n1678_40),
    .I2(u_usb_device_controller_usb_control_inst_s_sendbyte_7_16),
    .I3(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s9 .INIT=16'h00FE;
  LUT4 \u_usb_device_controller/u_usb_packet/s_state_11_s15  (
    .F(u_usb_device_controller_u_usb_packet_s_state_11),
    .I0(u_usb_device_controller_u_usb_packet_s_state_11_21),
    .I1(u_usb_device_controller_u_usb_packet_s_state_11_22),
    .I2(u_usb_device_controller_u_usb_packet_n624_37),
    .I3(u_usb_device_controller_u_usb_packet_s_state_11_23) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_11_s15 .INIT=16'h0B00;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s6  (
    .F(u_usb_device_controller_usb_transact_inst_s_sendpid_3_11),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3_13),
    .I1(u_usb_device_controller_usb_transact_inst_n1159_25),
    .I2(u_usb_device_controller_usb_transact_inst_s_in),
    .I3(u_usb_device_controller_usb_transact_inst_s_sendpid_3_14) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s6 .INIT=16'h0010;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1068_s6  (
    .F(u_usb_device_controller_usb_transact_inst_n1068_10),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I2(u_usb_device_controller_usb_transact_inst_n1111_22) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1068_s6 .INIT=8'h80;
  LUT4 \u_usb_device_controller/u_usb_packet/n640_s13  (
    .F(u_usb_device_controller_u_usb_packet_n640_18),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[3]),
    .I2(u_usb_device_controller_u_usb_packet_n640_27),
    .I3(u_usb_device_controller_u_usb_packet_n640_21) 
);
defparam \u_usb_device_controller/u_usb_packet/n640_s13 .INIT=16'h000B;
  LUT4 \u_usb_device_controller/u_usb_packet/n640_s14  (
    .F(u_usb_device_controller_u_usb_packet_n640_19),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[0]),
    .I1(u_usb_device_controller_u_usb_packet_n620),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf[8]),
    .I3(u_usb_device_controller_u_usb_packet_n622) 
);
defparam \u_usb_device_controller/u_usb_packet/n640_s14 .INIT=16'hB0BB;
  LUT4 \u_usb_device_controller/u_usb_packet/n642_s13  (
    .F(u_usb_device_controller_u_usb_packet_n642_18),
    .I0(u_usb_device_controller_u_usb_packet_n784_18),
    .I1(u_usb_device_controller_u_usb_packet_n782_8),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout[6]),
    .I3(u_usb_device_controller_u_usb_packet_n640_27) 
);
defparam \u_usb_device_controller/u_usb_packet/n642_s13 .INIT=16'h1F00;
  LUT4 \u_usb_device_controller/u_usb_packet/n642_s14  (
    .F(u_usb_device_controller_u_usb_packet_n642_19),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[2]),
    .I2(u_usb_device_controller_u_usb_packet_n642_21),
    .I3(u_usb_device_controller_u_usb_packet_n782_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n642_s14 .INIT=16'hF400;
  LUT4 \u_usb_device_controller/u_usb_packet/n642_s15  (
    .F(u_usb_device_controller_u_usb_packet_n642_20),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[1]),
    .I1(u_usb_device_controller_u_usb_packet_n620),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf[9]),
    .I3(u_usb_device_controller_u_usb_packet_n622) 
);
defparam \u_usb_device_controller/u_usb_packet/n642_s15 .INIT=16'hB0BB;
  LUT4 \u_usb_device_controller/u_usb_packet/n644_s13  (
    .F(u_usb_device_controller_u_usb_packet_n644_18),
    .I0(u_usb_device_controller_u_usb_packet_n784_18),
    .I1(u_usb_device_controller_u_usb_packet_n782_8),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout[5]),
    .I3(u_usb_device_controller_u_usb_packet_n640_27) 
);
defparam \u_usb_device_controller/u_usb_packet/n644_s13 .INIT=16'h1F00;
  LUT4 \u_usb_device_controller/u_usb_packet/n644_s14  (
    .F(u_usb_device_controller_u_usb_packet_n644_19),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[1]),
    .I2(u_usb_device_controller_u_usb_packet_n644_21),
    .I3(u_usb_device_controller_u_usb_packet_n782_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n644_s14 .INIT=16'hF400;
  LUT4 \u_usb_device_controller/u_usb_packet/n644_s15  (
    .F(u_usb_device_controller_u_usb_packet_n644_20),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[2]),
    .I1(u_usb_device_controller_u_usb_packet_n620),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf[10]),
    .I3(u_usb_device_controller_u_usb_packet_n622) 
);
defparam \u_usb_device_controller/u_usb_packet/n644_s15 .INIT=16'hB0BB;
  LUT4 \u_usb_device_controller/u_usb_packet/n646_s13  (
    .F(u_usb_device_controller_u_usb_packet_n646_18),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[0]),
    .I2(u_usb_device_controller_u_usb_packet_n640_27),
    .I3(u_usb_device_controller_u_usb_packet_n646_20) 
);
defparam \u_usb_device_controller/u_usb_packet/n646_s13 .INIT=16'h000B;
  LUT4 \u_usb_device_controller/u_usb_packet/n646_s14  (
    .F(u_usb_device_controller_u_usb_packet_n646_19),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[3]),
    .I1(u_usb_device_controller_u_usb_packet_n620),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf[11]),
    .I3(u_usb_device_controller_u_usb_packet_n622) 
);
defparam \u_usb_device_controller/u_usb_packet/n646_s14 .INIT=16'hB0BB;
  LUT3 \u_usb_device_controller/u_usb_packet/n650_s13  (
    .F(u_usb_device_controller_u_usb_packet_n650_18),
    .I0(u_usb_device_controller_u_usb_packet_n640_27),
    .I1(u_usb_device_controller_u_usb_packet_n650_20),
    .I2(u_usb_device_controller_u_usb_packet_n650_21) 
);
defparam \u_usb_device_controller/u_usb_packet/n650_s13 .INIT=8'h10;
  LUT4 \u_usb_device_controller/u_usb_packet/n650_s14  (
    .F(u_usb_device_controller_u_usb_packet_n650_19),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[5]),
    .I1(u_usb_device_controller_u_usb_packet_n620),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf[13]),
    .I3(u_usb_device_controller_u_usb_packet_n622) 
);
defparam \u_usb_device_controller/u_usb_packet/n650_s14 .INIT=16'hB0BB;
  LUT2 \u_usb_device_controller/u_usb_packet/n652_s13  (
    .F(u_usb_device_controller_u_usb_packet_n652_18),
    .I0(u_usb_device_controller_u_usb_packet_s_dataout[1]),
    .I1(u_usb_device_controller_u_usb_packet_n782_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n652_s13 .INIT=4'h8;
  LUT4 \u_usb_device_controller/u_usb_packet/n654_s13  (
    .F(u_usb_device_controller_u_usb_packet_n654_18),
    .I0(u_usb_device_controller_u_usb_packet_n626),
    .I1(u_usb_device_controller_u_usb_packet_n328_11),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout[0]),
    .I3(u_usb_device_controller_u_usb_packet_n782_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n654_s13 .INIT=16'h0777;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1064_s13  (
    .F(u_usb_device_controller_usb_transact_inst_n1064_18),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I1(u_usb_device_controller_usb_transact_inst_n1070_14),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1064_s13 .INIT=8'h10;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1066_s10  (
    .F(u_usb_device_controller_usb_transact_inst_n1066_14),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1066_s10 .INIT=4'h1;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1111_s14  (
    .F(u_usb_device_controller_usb_transact_inst_n1111_18),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1111_s14 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1074_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1074_23),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I2(u_usb_device_controller_usb_transact_inst_n1064_21),
    .I3(u_usb_device_controller_usb_transact_inst_s_in_valid) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1074_s18 .INIT=16'h4F00;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1074_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1074_24),
    .I0(u_usb_device_controller_usb_transact_inst_s_out),
    .I1(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I2(u_usb_device_controller_usb_transact_inst_s_in),
    .I3(u_usb_device_controller_usb_transact_inst_n1095_46) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1074_s19 .INIT=16'h0B33;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1070_s10  (
    .F(u_usb_device_controller_usb_transact_inst_n1070_14),
    .I0(u_usb_device_controller_usb_transact_inst_n1064_16),
    .I1(u_usb_device_controller_usb_transact_inst_n1064_27),
    .I2(u_usb_device_controller_usb_transact_inst_n1565_4),
    .I3(u_usb_device_controller_usb_transact_inst_n1070_20) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1070_s10 .INIT=16'h001F;
  LUT2 \u_usb_device_controller/usb_control_inst/n1672_s37  (
    .F(u_usb_device_controller_usb_control_inst_n1672_41),
    .I0(u_usb_device_controller_usb_control_inst_n1474_3),
    .I1(u_usb_device_controller_usb_control_inst_n1483_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s37 .INIT=4'h8;
  LUT4 \u_usb_device_controller/usb_control_inst/n1672_s38  (
    .F(u_usb_device_controller_usb_control_inst_n1672_42),
    .I0(u_usb_device_controller_usbc_dsclen_0_28),
    .I1(u_usb_device_controller_usb_control_inst_n1672_45),
    .I2(u_usb_device_controller_usb_control_inst_n1672_44),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscrd_4) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s38 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1672_s39  (
    .F(u_usb_device_controller_usb_control_inst_n1672_43),
    .I0(u_usb_device_controller_usb_transact_inst_txpop_o_d_9),
    .I1(u_usb_device_controller_usb_control_inst_n1672_46),
    .I2(u_usb_device_controller_usb_transact_inst_txpop_o_d_5),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_7_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s39 .INIT=16'h00EF;
  LUT3 \u_usb_device_controller/usb_control_inst/n1672_s40  (
    .F(u_usb_device_controller_usb_control_inst_n1672_44),
    .I0(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I1(u_usb_device_controller_u_usb_packet_n328_17),
    .I2(u_usb_device_controller_usb_transact_inst_s_in_valid) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s40 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1674_s35  (
    .F(u_usb_device_controller_usb_control_inst_n1674_39),
    .I0(u_usb_device_controller_usb_control_inst_n1674_44),
    .I1(u_usb_device_controller_usb_transact_inst_txpop_o_d_9),
    .I2(u_usb_device_controller_usb_control_inst_n1661_17),
    .I3(u_usb_device_controller_usb_control_inst_n1672_44) 
);
defparam \u_usb_device_controller/usb_control_inst/n1674_s35 .INIT=16'hD000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1676_s35  (
    .F(u_usb_device_controller_usb_control_inst_n1676_39),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]),
    .I3(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1676_s35 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/usb_control_inst/n1678_s36  (
    .F(u_usb_device_controller_usb_control_inst_n1678_40),
    .I0(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerptr_5_14) 
);
defparam \u_usb_device_controller/usb_control_inst/n1678_s36 .INIT=4'h8;
  LUT4 \u_usb_device_controller/usb_control_inst/n1678_s37  (
    .F(u_usb_device_controller_usb_control_inst_n1678_41),
    .I0(u_usb_device_controller_usb_control_inst_n1682_39),
    .I1(u_usb_device_controller_usb_control_inst_s_answerptr_5_10),
    .I2(u_usb_device_controller_usb_control_inst_n1678_43),
    .I3(u_usb_device_controller_usb_control_inst_n1678_44) 
);
defparam \u_usb_device_controller/usb_control_inst/n1678_s37 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1680_s38  (
    .F(u_usb_device_controller_usb_control_inst_n1680_42),
    .I0(u_usb_device_controller_usb_control_inst_n1680_50),
    .I1(u_usb_device_controller_usb_control_inst_n1670_39),
    .I2(u_usb_device_controller_usb_control_inst_n1680_46),
    .I3(u_usb_device_controller_usb_control_inst_n1629) 
);
defparam \u_usb_device_controller/usb_control_inst/n1680_s38 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/usb_control_inst/n1680_s39  (
    .F(u_usb_device_controller_usb_control_inst_n1680_43),
    .I0(u_usb_device_controller_usb_control_inst_n1680_47),
    .I1(u_usb_device_controller_usb_control_inst_n1672_44),
    .I2(u_usb_device_controller_usb_control_inst_n1682_39),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_5_10) 
);
defparam \u_usb_device_controller/usb_control_inst/n1680_s39 .INIT=16'h0700;
  LUT4 \u_usb_device_controller/usb_control_inst/n1680_s40  (
    .F(u_usb_device_controller_usb_control_inst_n1680_44),
    .I0(u_usb_device_controller_usb_control_inst_n1678_40),
    .I1(u_usb_device_controller_usb_control_inst_n1649_18),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_13),
    .I3(u_usb_device_controller_usb_control_inst_n1672_44) 
);
defparam \u_usb_device_controller/usb_control_inst/n1680_s40 .INIT=16'h00FE;
  LUT3 \u_usb_device_controller/usb_control_inst/n1682_s35  (
    .F(u_usb_device_controller_usb_control_inst_n1682_39),
    .I0(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I1(u_usb_device_controller_u_usb_packet_n328_17),
    .I2(u_usb_device_controller_usb_transact_inst_s_setup_2) 
);
defparam \u_usb_device_controller/usb_control_inst/n1682_s35 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1682_s36  (
    .F(u_usb_device_controller_usb_control_inst_n1682_40),
    .I0(u_usb_device_controller_usb_control_inst_n1836_15),
    .I1(u_usb_device_controller_usb_control_inst_n2067_7),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I3(u_usb_device_controller_usb_control_inst_s_interface_set_9) 
);
defparam \u_usb_device_controller/usb_control_inst/n1682_s36 .INIT=16'h007F;
  LUT3 \u_usb_device_controller/usb_control_inst/n1684_s35  (
    .F(u_usb_device_controller_usb_control_inst_n1684_39),
    .I0(u_usb_device_controller_usb_control_inst_s_state[2]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[3]),
    .I2(u_usb_device_controller_usb_control_inst_n1684_41) 
);
defparam \u_usb_device_controller/usb_control_inst/n1684_s35 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1684_s36  (
    .F(u_usb_device_controller_usb_control_inst_n1684_40),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I3(u_usb_device_controller_usb_control_inst_n1684_42) 
);
defparam \u_usb_device_controller/usb_control_inst/n1684_s36 .INIT=16'h0001;
  LUT3 \u_usb_device_controller/usb_control_inst/n1686_s35  (
    .F(u_usb_device_controller_usb_control_inst_n1686_39),
    .I0(u_usb_device_controller_usb_control_inst_s_state[3]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[2]),
    .I2(u_usb_device_controller_usb_control_inst_n1684_41) 
);
defparam \u_usb_device_controller/usb_control_inst/n1686_s35 .INIT=8'h40;
  LUT3 \u_usb_device_controller/usb_control_inst/n1686_s36  (
    .F(u_usb_device_controller_usb_control_inst_n1686_40),
    .I0(u_usb_device_controller_usb_control_inst_n1836_15),
    .I1(u_usb_device_controller_usb_control_inst_n1686_41),
    .I2(u_usb_device_controller_usb_control_inst_n1686_42) 
);
defparam \u_usb_device_controller/usb_control_inst/n1686_s36 .INIT=8'h20;
  LUT4 \u_usb_device_controller/usb_control_inst/n1688_s35  (
    .F(u_usb_device_controller_usb_control_inst_n1688_39),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I1(u_usb_device_controller_usb_control_inst_n1682_39),
    .I2(u_usb_device_controller_usb_control_inst_n1686_41),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/usb_control_inst/n1688_s35 .INIT=16'h0FBB;
  LUT4 \u_usb_device_controller/usb_control_inst/n1690_s30  (
    .F(u_usb_device_controller_usb_control_inst_n1690_34),
    .I0(u_usb_device_controller_usb_control_inst_s_answerptr_7_12),
    .I1(u_usb_device_controller_n2393_9),
    .I2(u_usb_device_controller_usb_control_inst_n1686_39),
    .I3(u_usb_device_controller_usb_control_inst_n1690_37) 
);
defparam \u_usb_device_controller/usb_control_inst/n1690_s30 .INIT=16'h000D;
  LUT4 \u_usb_device_controller/usb_control_inst/n1690_s31  (
    .F(u_usb_device_controller_usb_control_inst_n1690_35),
    .I0(u_usb_device_controller_usb_control_inst_n2896_9),
    .I1(u_usb_device_controller_usb_control_inst_n1690_38),
    .I2(u_usb_device_controller_usb_control_inst_n1670_43),
    .I3(u_usb_device_controller_usb_control_inst_n1682_39) 
);
defparam \u_usb_device_controller/usb_control_inst/n1690_s31 .INIT=16'h00F8;
  LUT4 \u_usb_device_controller/usb_control_inst/n1690_s32  (
    .F(u_usb_device_controller_usb_control_inst_n1690_36),
    .I0(u_usb_device_controller_usb_control_inst_n1672_45),
    .I1(u_usb_device_controller_usbc_dsclen_0_28),
    .I2(u_usb_device_controller_usb_control_inst_n1672_44),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscrd_4) 
);
defparam \u_usb_device_controller/usb_control_inst/n1690_s32 .INIT=16'hE000;
  LUT3 \u_usb_device_controller/usb_control_inst/n1701_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1701_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1701_s12 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_control_inst/n1701_s13  (
    .F(u_usb_device_controller_usb_control_inst_n1701_17),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I2(u_usb_device_controller_usb_control_inst_n1701_21) 
);
defparam \u_usb_device_controller/usb_control_inst/n1701_s13 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1701_s14  (
    .F(u_usb_device_controller_usb_control_inst_n1701_18),
    .I0(u_usb_device_controller_usb_control_inst_n1876_9),
    .I1(u_usb_device_controller_usb_control_inst_n1701_21),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1876_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1701_s14 .INIT=16'h8F00;
  LUT3 \u_usb_device_controller/usb_control_inst/n1703_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1703_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1703_s12 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_control_inst/n1705_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1705_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1705_s12 .INIT=8'h40;
  LUT3 \u_usb_device_controller/usb_control_inst/n1707_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1707_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1707_s12 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_control_inst/n1711_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1711_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1711_s12 .INIT=8'h40;
  LUT3 \u_usb_device_controller/usb_control_inst/n1713_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1713_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1713_s12 .INIT=8'h80;
  LUT3 \u_usb_device_controller/usb_control_inst/n1715_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1715_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1715_s12 .INIT=8'h01;
  LUT3 \u_usb_device_controller/usb_control_inst/n1715_s13  (
    .F(u_usb_device_controller_usb_control_inst_n1715_17),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I2(u_usb_device_controller_usb_control_inst_n1701_21) 
);
defparam \u_usb_device_controller/usb_control_inst/n1715_s13 .INIT=8'h80;
  LUT3 \u_usb_device_controller/usb_control_inst/n1731_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1731_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I2(u_usb_device_controller_usb_control_inst_n1701_21) 
);
defparam \u_usb_device_controller/usb_control_inst/n1731_s12 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_control_inst/n1745_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1745_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_n1701_21) 
);
defparam \u_usb_device_controller/usb_control_inst/n1745_s12 .INIT=8'h40;
  LUT3 \u_usb_device_controller/usb_control_inst/n1775_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1775_13),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I2(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1775_s9 .INIT=8'h80;
  LUT3 \u_usb_device_controller/usb_control_inst/n1805_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1805_13),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1805_s9 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1649_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1649_16),
    .I0(u_usb_device_controller_usb_control_inst_s_sendbyte_7_15),
    .I1(u_usb_device_controller_usb_control_inst_n1649_19),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscoff[5]),
    .I3(u_usb_device_controller_usb_control_inst_n1678_40) 
);
defparam \u_usb_device_controller/usb_control_inst/n1649_s12 .INIT=16'h7800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1649_s13  (
    .F(u_usb_device_controller_usb_control_inst_n1649_17),
    .I0(u_usb_device_controller_usb_control_inst_s_sendbyte_7_15),
    .I1(u_usb_device_controller_usb_control_inst_n1649_23),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscrd_4),
    .I3(u_usb_device_controller_usb_control_inst_n1649_19) 
);
defparam \u_usb_device_controller/usb_control_inst/n1649_s13 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_control_inst/n1649_s14  (
    .F(u_usb_device_controller_usb_control_inst_n1649_18),
    .I0(u_usb_device_controller_usb_control_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[5]),
    .I2(u_usb_device_controller_usb_control_inst_n1629_4),
    .I3(u_usb_device_controller_usb_control_inst_n1649_21) 
);
defparam \u_usb_device_controller/usb_control_inst/n1649_s14 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1652_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1652_16),
    .I0(u_usb_device_controller_usb_control_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[5]),
    .I2(u_usb_device_controller_usb_control_inst_n1629_4),
    .I3(u_usb_device_controller_usb_control_inst_n1652_19) 
);
defparam \u_usb_device_controller/usb_control_inst/n1652_s12 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/usb_control_inst/n1652_s14  (
    .F(u_usb_device_controller_usb_control_inst_n1652_18),
    .I0(u_usb_device_controller_usb_control_inst_n1652_22),
    .I1(u_usb_device_controller_usb_control_inst_s_sendbyte_7_15),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscrd_4) 
);
defparam \u_usb_device_controller/usb_control_inst/n1652_s14 .INIT=8'h0B;
  LUT2 \u_usb_device_controller/usb_control_inst/n1658_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1658_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1658_s12 .INIT=4'h8;
  LUT4 \u_usb_device_controller/usb_control_inst/n1661_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1661_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_sendbyte_7_15),
    .I2(u_usb_device_controller_usb_control_inst_n1672_41),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1661_s12 .INIT=16'h7F80;
  LUT4 \u_usb_device_controller/usb_control_inst/n1661_s13  (
    .F(u_usb_device_controller_usb_control_inst_n1661_17),
    .I0(u_usb_device_controller_usb_control_inst_s_state[7]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[8]),
    .I3(u_usb_device_controller_usb_control_inst_n1661_22) 
);
defparam \u_usb_device_controller/usb_control_inst/n1661_s13 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1661_s14  (
    .F(u_usb_device_controller_usb_control_inst_n1661_18),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_sendbyte_7_15),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]),
    .I3(u_usb_device_controller_usb_control_inst_n1678_40) 
);
defparam \u_usb_device_controller/usb_control_inst/n1661_s14 .INIT=16'h7800;
  LUT3 \u_usb_device_controller/usb_control_inst/n1661_s15  (
    .F(u_usb_device_controller_usb_control_inst_n1661_19),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscrd_4) 
);
defparam \u_usb_device_controller/usb_control_inst/n1661_s15 .INIT=8'h60;
  LUT3 \u_usb_device_controller/u_usb_packet/n620_s42  (
    .F(u_usb_device_controller_u_usb_packet_n620_47),
    .I0(u_usb_device_controller_u_usb_packet_s_state[8]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[7]),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout_7_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n620_s42 .INIT=8'h40;
  LUT3 \u_usb_device_controller/u_usb_packet/n626_s37  (
    .F(u_usb_device_controller_u_usb_packet_n626_41),
    .I0(u_usb_device_controller_usb_transact_inst_n1080_53),
    .I1(u_usb_device_controller_usb_transact_inst_n1072_18),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_28) 
);
defparam \u_usb_device_controller/u_usb_packet/n626_s37 .INIT=8'h9B;
  LUT4 \u_usb_device_controller/u_usb_packet/n626_s38  (
    .F(u_usb_device_controller_u_usb_packet_n626_42),
    .I0(u_usb_device_controller_u_usb_packet_n626_44),
    .I1(u_usb_device_controller_usb_control_inst_n1652_16),
    .I2(u_usb_device_controller_u_usb_packet_n626_45),
    .I3(u_usb_device_controller_usb_transact_inst_txpop_o_d_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n626_s38 .INIT=16'h0D00;
  LUT4 \u_usb_device_controller/u_usb_packet/n628_s43  (
    .F(u_usb_device_controller_u_usb_packet_n628_47),
    .I0(u_usb_device_controller_u_usb_packet_s_rxerror),
    .I1(u_usb_device_controller_usb_transact_inst_n1565_4),
    .I2(u_usb_device_controller_u_usb_packet_s_state_11_22),
    .I3(u_usb_device_controller_u_usb_packet_n628_48) 
);
defparam \u_usb_device_controller/u_usb_packet/n628_s43 .INIT=16'h4000;
  LUT3 \u_usb_device_controller/u_usb_packet/n633_s35  (
    .F(u_usb_device_controller_u_usb_packet_n633_39),
    .I0(u_usb_device_controller_u_usb_packet_n633_40),
    .I1(u_usb_device_controller_u_usb_packet_n633_41),
    .I2(u_usb_device_controller_u_usb_packet_n633_42) 
);
defparam \u_usb_device_controller/u_usb_packet/n633_s35 .INIT=8'h01;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1088_s40  (
    .F(u_usb_device_controller_usb_transact_inst_n1088_44),
    .I0(u_usb_device_controller_usb_transact_inst_n1088_48),
    .I1(u_usb_device_controller_usb_transact_inst_n1086_48) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1088_s40 .INIT=4'h1;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1088_s41  (
    .F(u_usb_device_controller_usb_transact_inst_n1088_45),
    .I0(u_usb_device_controller_u_usb_packet_n626_42),
    .I1(u_usb_device_controller_usb_transact_inst_txpop_o_d_5),
    .I2(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_24) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1088_s41 .INIT=16'hF0BB;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1090_s42  (
    .F(u_usb_device_controller_usb_transact_inst_n1090_46),
    .I0(u_usb_device_controller_usb_transact_inst_s_prevrxact),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I2(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I3(u_usb_device_controller_usb_transact_inst_n1105_48) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1090_s42 .INIT=16'h00FE;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1091_s44  (
    .F(u_usb_device_controller_usb_transact_inst_n1091_49),
    .I0(u_usb_device_controller_usb_transact_inst_n1091_54),
    .I1(u_usb_device_controller_u_usb_packet_n800_6) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1091_s44 .INIT=4'h1;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1091_s45  (
    .F(u_usb_device_controller_usb_transact_inst_n1091_50),
    .I0(u_usb_device_controller_usb_transact_inst_n1157_27),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_28),
    .I2(u_usb_device_controller_usb_transact_inst_n1041_4),
    .I3(u_usb_device_controller_usb_transact_inst_n1091_52) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1091_s45 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1093_s47  (
    .F(u_usb_device_controller_usb_transact_inst_n1093_51),
    .I0(u_usb_device_controller_usb_transact_inst_n1080_55),
    .I1(u_usb_device_controller_usb_transact_inst_n1105_48),
    .I2(u_usb_device_controller_u_usb_packet_n626_41),
    .I3(u_usb_device_controller_usb_transact_inst_n1091_49) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1093_s47 .INIT=16'hB0BB;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1095_s40  (
    .F(u_usb_device_controller_usb_transact_inst_n1095_44),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1095_s40 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1095_s41  (
    .F(u_usb_device_controller_usb_transact_inst_n1095_45),
    .I0(u_usb_device_controller_usb_transact_inst_n1157_26),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_27),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_28),
    .I3(u_usb_device_controller_usb_transact_inst_n1095_47) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1095_s41 .INIT=16'h8000;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1095_s42  (
    .F(u_usb_device_controller_usb_transact_inst_n1095_46),
    .I0(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I1(u_usb_device_controller_u_usb_packet_s_rxerror),
    .I2(u_usb_device_controller_u_usb_packet_s_rxgoodpacket) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1095_s42 .INIT=8'h10;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1099_s43  (
    .F(u_usb_device_controller_usb_transact_inst_n1099_47),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3_11),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid_3_21),
    .I2(u_usb_device_controller_usb_transact_inst_n1093_51),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[5]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1099_s43 .INIT=16'hB0BB;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1101_s40  (
    .F(u_usb_device_controller_usb_transact_inst_n1101_44),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3_11),
    .I1(u_usb_device_controller_usb_transact_inst_n1101_45),
    .I2(u_usb_device_controller_usb_transact_inst_n1105_48),
    .I3(u_usb_device_controller_usb_transact_inst_n1101_48) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1101_s40 .INIT=16'hFE00;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1105_s43  (
    .F(u_usb_device_controller_usb_transact_inst_n1105_47),
    .I0(u_usb_device_controller_usb_transact_inst_s_sof),
    .I1(u_usb_device_controller_usb_transact_inst_n1159_25),
    .I2(u_usb_device_controller_usb_transact_inst_n162_3) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1105_s43 .INIT=8'h10;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1105_s44  (
    .F(u_usb_device_controller_usb_transact_inst_n1105_48),
    .I0(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1105_s44 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1109_s43  (
    .F(u_usb_device_controller_usb_transact_inst_n1109_47),
    .I0(u_usb_device_controller_usb_transact_inst_n1064_27),
    .I1(u_usb_device_controller_usb_transact_inst_n1109_49),
    .I2(u_usb_device_controller_usb_transact_inst_n1080),
    .I3(u_usb_device_controller_u_usb_packet_usbp_rxact) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1109_s43 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1109_s44  (
    .F(u_usb_device_controller_usb_transact_inst_n1109_48),
    .I0(u_usb_device_controller_usb_transact_inst_n1088_48),
    .I1(u_usb_device_controller_usb_transact_inst_n1070_20),
    .I2(u_usb_device_controller_usb_transact_inst_s_endpt_0_9),
    .I3(u_usb_device_controller_usb_transact_inst_n1105_47) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1109_s44 .INIT=16'h0BBB;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1138_s24  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_29),
    .I0(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I1(u_usb_device_controller_usb_transact_inst_n1142_25) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s24 .INIT=4'h1;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1138_s25  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_30),
    .I0(u_usb_device_controller_usb_transact_inst_n1138_35),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[7]),
    .I2(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[8]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s25 .INIT=16'h0D00;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1140_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1140_22),
    .I0(u_usb_device_controller_usb_transact_inst_n1138_37),
    .I1(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I2(u_usb_device_controller_usb_transact_inst_wait_count[7]),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_35) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1140_s18 .INIT=16'h0130;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1142_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1142_23),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[4]),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[5]),
    .I2(u_usb_device_controller_usb_transact_inst_n1146_22) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1142_s19 .INIT=8'h10;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1144_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1144_22),
    .I0(u_usb_device_controller_usb_transact_inst_n1146_22),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[4]),
    .I2(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[5]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1144_s18 .INIT=16'h0D00;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1146_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1146_22),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[0]),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[1]),
    .I2(u_usb_device_controller_usb_transact_inst_wait_count[2]),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[3]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1146_s18 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1148_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1148_22),
    .I0(u_usb_device_controller_usb_transact_inst_n1150_22),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[2]),
    .I2(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[3]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1148_s18 .INIT=16'h0D00;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1150_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1150_22),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[0]),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[1]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1150_s18 .INIT=4'h1;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1152_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1152_22),
    .I0(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[1]),
    .I2(u_usb_device_controller_usb_transact_inst_wait_count[0]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1152_s18 .INIT=8'h40;
  LUT4 \u_usb_device_controller/n1615_s10  (
    .F(u_usb_device_controller_n1615_15),
    .I0(u_usb_device_controller_cur_state[0]),
    .I1(u_usb_device_controller_cur_state[1]),
    .I2(u_usb_device_controller_cur_state[3]),
    .I3(u_usb_device_controller_cur_state[2]) 
);
defparam \u_usb_device_controller/n1615_s10 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1076_s15  (
    .F(u_usb_device_controller_usb_transact_inst_n1076_21),
    .I0(u_usb_device_controller_usb_transact_inst_s_out),
    .I1(u_usb_device_controller_usb_transact_inst_s_out_valid),
    .I2(u_usb_device_controller_usb_transact_inst_s_in),
    .I3(u_usb_device_controller_usb_transact_inst_n1095_46) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1076_s15 .INIT=16'h0ECC;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1072_s14  (
    .F(u_usb_device_controller_usb_transact_inst_n1072_20),
    .I0(u_usb_device_controller_usb_transact_inst_n1072_22),
    .I1(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I2(u_usb_device_controller_usb_transact_inst_n1072_18),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[5]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1072_s14 .INIT=16'hD000;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1157_s24  (
    .F(u_usb_device_controller_usb_transact_inst_n1157_30),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[6]),
    .I1(u_usb_device_controller_s_isync),
    .I2(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1157_s24 .INIT=8'hA3;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1157_s25  (
    .F(u_usb_device_controller_usb_transact_inst_n1157_31),
    .I0(u_usb_device_controller_usb_transact_inst_n1159_25),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid_3_13),
    .I2(u_usb_device_controller_usb_transact_inst_s_sendpid_3_14),
    .I3(u_usb_device_controller_usb_transact_inst_s_sendpid_3_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1157_s25 .INIT=16'h00FE;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1159_s20  (
    .F(u_usb_device_controller_usb_transact_inst_n1159_25),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_test_en),
    .I2(u_usb_device_controller_utmi_dataout_o_d_0_4) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1159_s20 .INIT=8'h80;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1159_s21  (
    .F(u_usb_device_controller_usb_transact_inst_n1159_26),
    .I0(u_usb_device_controller_usb_transact_inst_n1159_27),
    .I1(u_usb_device_controller_usb_transact_inst_n1099_49),
    .I2(u_usb_device_controller_usb_transact_inst_s_sendpid_3_14) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1159_s21 .INIT=8'h07;
  LUT3 \u_usb_device_controller/usb_control_inst/n1860_s24  (
    .F(u_usb_device_controller_usb_control_inst_n1860_29),
    .I0(u_usb_device_controller_usb_control_inst_n1860_31),
    .I1(u_usb_device_controller_usb_control_inst_n645_51),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1860_s24 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/usb_control_inst/n1860_s25  (
    .F(u_usb_device_controller_usb_control_inst_n1860_30),
    .I0(u_usb_device_controller_usb_control_inst_n1860_32),
    .I1(u_usb_device_controller_usb_control_inst_usbc_txdat[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_sendbyte_7_14),
    .I3(u_usb_device_controller_usb_control_inst_n2896_4) 
);
defparam \u_usb_device_controller/usb_control_inst/n1860_s25 .INIT=16'hAC00;
  LUT4 \u_usb_device_controller/n385_s3  (
    .F(u_usb_device_controller_n385_7),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I2(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I3(u_usb_device_controller_rxact_o_d) 
);
defparam \u_usb_device_controller/n385_s3 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/n443_s3  (
    .F(u_usb_device_controller_n443_7),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .I2(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I3(u_usb_device_controller_rxact_o_d) 
);
defparam \u_usb_device_controller/n443_s3 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/n503_s3  (
    .F(u_usb_device_controller_n503_7),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .I2(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I3(u_usb_device_controller_rxact_o_d) 
);
defparam \u_usb_device_controller/n503_s3 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/n561_s3  (
    .F(u_usb_device_controller_n561_7),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .I2(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I3(u_usb_device_controller_rxact_o_d) 
);
defparam \u_usb_device_controller/n561_s3 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/s_ctlparam_7_s4  (
    .F(u_usb_device_controller_usb_control_inst_s_ctlparam_7_7),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I1(u_usb_device_controller_usb_control_inst_n1864_8),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .I3(u_usb_device_controller_usb_control_inst_s_ctlparam_7_8) 
);
defparam \u_usb_device_controller/usb_control_inst/s_ctlparam_7_s4 .INIT=16'h001F;
  LUT3 \u_usb_device_controller/isync_1_s5  (
    .F(u_usb_device_controller_isync_1_10),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I2(u_usb_device_controller_txpktfin_o_d) 
);
defparam \u_usb_device_controller/isync_1_s5 .INIT=8'h40;
  LUT3 \u_usb_device_controller/isync_2_s4  (
    .F(u_usb_device_controller_isync_2_9),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .I2(u_usb_device_controller_txpktfin_o_d) 
);
defparam \u_usb_device_controller/isync_2_s4 .INIT=8'h40;
  LUT3 \u_usb_device_controller/isync_3_s4  (
    .F(u_usb_device_controller_isync_3_9),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .I2(u_usb_device_controller_txpktfin_o_d) 
);
defparam \u_usb_device_controller/isync_3_s4 .INIT=8'h80;
  LUT3 \u_usb_device_controller/isync_4_s5  (
    .F(u_usb_device_controller_isync_4_10),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .I2(u_usb_device_controller_txpktfin_o_d) 
);
defparam \u_usb_device_controller/isync_4_s5 .INIT=8'h10;
  LUT4 \u_usb_device_controller/test_packet_inst/cnt_11_s4  (
    .F(u_usb_device_controller_test_packet_inst_cnt_11_9),
    .I0(u_usb_device_controller_test_packet_inst_n133_6),
    .I1(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I2(u_usb_device_controller_test_packet_inst_cnt_11_11),
    .I3(u_usb_device_controller_test_packet_inst_n318_9) 
);
defparam \u_usb_device_controller/test_packet_inst/cnt_11_s4 .INIT=16'h1F00;
  LUT3 \u_usb_device_controller/test_packet_inst/cnt_11_s5  (
    .F(u_usb_device_controller_test_packet_inst_cnt_11_10),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_test_packet_inst_cnt_11_12),
    .I2(u_usb_device_controller_test_packet_inst_cnt_11_13) 
);
defparam \u_usb_device_controller/test_packet_inst/cnt_11_s5 .INIT=8'h40;
  LUT4 \u_usb_device_controller/test_packet_inst/test_data_6_s4  (
    .F(u_usb_device_controller_test_packet_inst_test_data_6),
    .I0(u_usb_device_controller_test_packet_inst_cnt[4]),
    .I1(u_usb_device_controller_test_packet_inst_test_data_6_9),
    .I2(u_usb_device_controller_test_packet_inst_cnt[5]),
    .I3(u_usb_device_controller_test_packet_inst_n318_9) 
);
defparam \u_usb_device_controller/test_packet_inst/test_data_6_s4 .INIT=16'h4F00;
  LUT4 \u_usb_device_controller/test_packet_inst/test_data_6_s5  (
    .F(u_usb_device_controller_test_packet_inst_test_data_6_8),
    .I0(u_usb_device_controller_test_packet_inst_cnt_11_9),
    .I1(u_usb_device_controller_test_packet_inst_n378_8),
    .I2(utmi_txready_i_d),
    .I3(u_usb_device_controller_test_packet_inst_test_en_dly_Z) 
);
defparam \u_usb_device_controller/test_packet_inst/test_data_6_s5 .INIT=16'h0700;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_2_s9  (
    .F(u_usb_device_controller_u_usb_init_s_state_2_14),
    .I0(u_usb_device_controller_u_usb_init_s_state[3]),
    .I1(u_usb_device_controller_u_usb_init_s_state_2_20),
    .I2(u_usb_device_controller_u_usb_init_n217_38),
    .I3(u_usb_device_controller_u_usb_init_s_state_2_16) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_2_s9 .INIT=16'h00EF;
  LUT4 \u_usb_device_controller/test_packet_inst/n318_s4  (
    .F(u_usb_device_controller_test_packet_inst_n318_8),
    .I0(u_usb_device_controller_test_packet_inst_n318_11),
    .I1(u_usb_device_controller_test_packet_inst_n133_7),
    .I2(u_usb_device_controller_test_packet_inst_n318_12),
    .I3(u_usb_device_controller_test_packet_inst_cnt[5]) 
);
defparam \u_usb_device_controller/test_packet_inst/n318_s4 .INIT=16'h0FBB;
  LUT3 \u_usb_device_controller/test_packet_inst/n318_s5  (
    .F(u_usb_device_controller_test_packet_inst_n318_9),
    .I0(u_usb_device_controller_test_packet_inst_cnt[6]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[7]),
    .I2(u_usb_device_controller_test_packet_inst_n318_13) 
);
defparam \u_usb_device_controller/test_packet_inst/n318_s5 .INIT=8'h10;
  LUT4 \u_usb_device_controller/test_packet_inst/n318_s6  (
    .F(u_usb_device_controller_test_packet_inst_n318_10),
    .I0(utmi_txready_i_d),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_test_packet_inst_n318_14),
    .I3(u_usb_device_controller_test_packet_inst_n318_17) 
);
defparam \u_usb_device_controller/test_packet_inst/n318_s6 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/test_packet_inst/n317_s5  (
    .F(u_usb_device_controller_test_packet_inst_n317_9),
    .I0(u_usb_device_controller_test_packet_inst_cnt_11_11),
    .I1(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I2(u_usb_device_controller_test_packet_inst_n318_9),
    .I3(u_usb_device_controller_test_packet_inst_n317_11) 
);
defparam \u_usb_device_controller/test_packet_inst/n317_s5 .INIT=16'h7000;
  LUT4 \u_usb_device_controller/test_packet_inst/n317_s6  (
    .F(u_usb_device_controller_test_packet_inst_n317_10),
    .I0(u_usb_device_controller_test_packet_inst_n314_8),
    .I1(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I2(u_usb_device_controller_test_packet_inst_n318_14),
    .I3(u_usb_device_controller_test_packet_inst_test_en_dly_Z) 
);
defparam \u_usb_device_controller/test_packet_inst/n317_s6 .INIT=16'h4F00;
  LUT4 \u_usb_device_controller/test_packet_inst/n312_s4  (
    .F(u_usb_device_controller_test_packet_inst_n312_8),
    .I0(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[2]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I3(u_usb_device_controller_test_packet_inst_test_data_val_9) 
);
defparam \u_usb_device_controller/test_packet_inst/n312_s4 .INIT=16'hBF00;
  LUT4 \u_usb_device_controller/test_packet_inst/n312_s5  (
    .F(u_usb_device_controller_test_packet_inst_n312_9),
    .I0(u_usb_device_controller_test_packet_inst_cnt_11_11),
    .I1(u_usb_device_controller_test_packet_inst_cnt_11_9),
    .I2(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I3(u_usb_device_controller_test_packet_inst_test_data_6) 
);
defparam \u_usb_device_controller/test_packet_inst/n312_s5 .INIT=16'h007F;
  LUT4 \u_usb_device_controller/test_packet_inst/n312_s6  (
    .F(u_usb_device_controller_test_packet_inst_n312_10),
    .I0(u_usb_device_controller_test_packet_inst_n318_17),
    .I1(u_usb_device_controller_test_packet_inst_cnt[4]),
    .I2(u_usb_device_controller_test_packet_inst_n312_13),
    .I3(u_usb_device_controller_test_packet_inst_test_en_dly_Z) 
);
defparam \u_usb_device_controller/test_packet_inst/n312_s6 .INIT=16'h4F00;
  LUT3 \u_usb_device_controller/test_packet_inst/n311_s5  (
    .F(u_usb_device_controller_test_packet_inst_n311_9),
    .I0(u_usb_device_controller_test_packet_inst_n311_10),
    .I1(u_usb_device_controller_test_packet_inst_cnt_11_9),
    .I2(u_usb_device_controller_test_packet_inst_test_data_6) 
);
defparam \u_usb_device_controller/test_packet_inst/n311_s5 .INIT=8'h0B;
  LUT4 \u_usb_device_controller/u_usb_init/n213_s20  (
    .F(u_usb_device_controller_u_usb_init_n213_28),
    .I0(u_usb_device_controller_u_usb_init_s_state[1]),
    .I1(u_usb_device_controller_u_usb_init_s_state[2]),
    .I2(u_usb_device_controller_u_usb_init_n212_57),
    .I3(u_usb_device_controller_u_usb_init_n212_39) 
);
defparam \u_usb_device_controller/u_usb_init/n213_s20 .INIT=16'h6000;
  LUT4 \u_usb_device_controller/u_usb_init/n219_s20  (
    .F(u_usb_device_controller_u_usb_init_n219_28),
    .I0(u_usb_device_controller_u_usb_init_n215_53),
    .I1(u_usb_device_controller_u_usb_init_s_state[1]),
    .I2(u_usb_device_controller_u_usb_init_s_state[2]),
    .I3(u_usb_device_controller_u_usb_init_n219_29) 
);
defparam \u_usb_device_controller/u_usb_init/n219_s20 .INIT=16'hD73F;
  LUT4 \u_usb_device_controller/n1534_s19  (
    .F(u_usb_device_controller_n1534_26),
    .I0(u_usb_device_controller_n1810_6),
    .I1(u_usb_device_controller_n2393_9),
    .I2(u_usb_device_controller_cur_state[0]),
    .I3(u_usb_device_controller_n1529_31) 
);
defparam \u_usb_device_controller/n1534_s19 .INIT=16'hB000;
  LUT4 \u_usb_device_controller/n1534_s21  (
    .F(u_usb_device_controller_n1534_28),
    .I0(u_usb_device_controller_usb_transact_inst_n1072_22),
    .I1(u_usb_device_controller_usb_transact_inst_txpop_o_d_5),
    .I2(u_usb_device_controller_n1473_50),
    .I3(u_usb_device_controller_cur_state[0]) 
);
defparam \u_usb_device_controller/n1534_s21 .INIT=16'h00BF;
  LUT4 \u_usb_device_controller/n1534_s22  (
    .F(u_usb_device_controller_n1534_29),
    .I0(u_usb_device_controller_n1534_32),
    .I1(u_usb_device_controller_n1534_33),
    .I2(u_usb_device_controller_n1534_34),
    .I3(u_usb_device_controller_n1529_25) 
);
defparam \u_usb_device_controller/n1534_s22 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/n1529_s18  (
    .F(u_usb_device_controller_n1529_24),
    .I0(u_usb_device_controller_s_halt_out),
    .I1(u_usb_device_controller_rxdat_d0_7_9),
    .I2(u_usb_device_controller_cur_state[1]),
    .I3(u_usb_device_controller_cur_state[0]) 
);
defparam \u_usb_device_controller/n1529_s18 .INIT=16'h00F4;
  LUT4 \u_usb_device_controller/n1529_s19  (
    .F(u_usb_device_controller_n1529_25),
    .I0(u_usb_device_controller_usb_transact_inst_T_PING_2),
    .I1(u_usb_device_controller_rxdat_d0_7_9),
    .I2(u_usb_device_controller_n1534_30),
    .I3(u_usb_device_controller_n1585_4) 
);
defparam \u_usb_device_controller/n1529_s19 .INIT=16'hFE00;
  LUT4 \u_usb_device_controller/n1529_s20  (
    .F(u_usb_device_controller_n1529_26),
    .I0(u_usb_device_controller_n1529_28),
    .I1(u_usb_device_controller_s_halt_in),
    .I2(u_usb_device_controller_n1534_30),
    .I3(u_usb_device_controller_n1529_29) 
);
defparam \u_usb_device_controller/n1529_s20 .INIT=16'h3A00;
  LUT4 \u_usb_device_controller/n1524_s19  (
    .F(u_usb_device_controller_n1524_25),
    .I0(u_usb_device_controller_n2393_9),
    .I1(u_usb_device_controller_n1810_6),
    .I2(u_usb_device_controller_cur_state[0]),
    .I3(u_usb_device_controller_n1529_31) 
);
defparam \u_usb_device_controller/n1524_s19 .INIT=16'hDF00;
  LUT3 \u_usb_device_controller/usbc_dsclen_0_s10  (
    .F(u_usb_device_controller_usbc_dsclen_0_15),
    .I0(u_usb_device_controller_usbc_dsclen_0_18),
    .I1(u_usb_device_controller_usbc_dsclen_0_19),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s10 .INIT=8'h35;
  LUT4 \u_usb_device_controller/usbc_dsclen_1_s9  (
    .F(u_usb_device_controller_usbc_dsclen_1_14),
    .I0(desc_qual_len_i_d[1]),
    .I1(u_usb_device_controller_usbc_dsclen_1_16),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s9 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/usbc_dsclen_1_s10  (
    .F(u_usb_device_controller_usbc_dsclen_1_15),
    .I0(u_usb_device_controller_usbc_dsclen_1_26),
    .I1(u_usb_device_controller_usbc_dsclen_1_18),
    .I2(u_usb_device_controller_usbc_dsclen_1_24),
    .I3(u_usb_device_controller_usbc_dsclen_1_20) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s10 .INIT=16'h4F00;
  LUT3 \u_usb_device_controller/usbc_dsclen_2_s9  (
    .F(u_usb_device_controller_usbc_dsclen_2_14),
    .I0(desc_dev_len_i_d[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_usbc_dsclen_2_16) 
);
defparam \u_usb_device_controller/usbc_dsclen_2_s9 .INIT=8'h0D;
  LUT4 \u_usb_device_controller/usbc_dsclen_2_s10  (
    .F(u_usb_device_controller_usbc_dsclen_2_15),
    .I0(u_usb_device_controller_usbc_dsclen_2_17),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_len_i_d[2]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/usbc_dsclen_2_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/usbc_dsclen_3_s9  (
    .F(u_usb_device_controller_usbc_dsclen_3_14),
    .I0(u_usb_device_controller_usbc_dsclen_3_15),
    .I1(u_usb_device_controller_usbc_dsclen_3_16),
    .I2(u_usb_device_controller_usbc_dsclen_3_17),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_3_s9 .INIT=16'h0FEE;
  LUT4 \u_usb_device_controller/usbc_dsclen_4_s9  (
    .F(u_usb_device_controller_usbc_dsclen_4_14),
    .I0(desc_dev_len_i_d[4]),
    .I1(u_usb_device_controller_usbc_dsclen_4_16),
    .I2(u_usb_device_controller_usbc_dsclen_4_17),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_4_s9 .INIT=16'h0305;
  LUT4 \u_usb_device_controller/usbc_dsclen_4_s10  (
    .F(u_usb_device_controller_usbc_dsclen_4_15),
    .I0(u_usb_device_controller_usbc_dsclen_4_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_len_i_d[4]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/usbc_dsclen_4_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/usbc_dsclen_5_s9  (
    .F(u_usb_device_controller_usbc_dsclen_5_14),
    .I0(u_usb_device_controller_usbc_dsclen_5_15),
    .I1(u_usb_device_controller_usbc_dsclen_5_16),
    .I2(u_usb_device_controller_usbc_dsclen_5_17),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_5_s9 .INIT=16'h0FBB;
  LUT2 \u_usb_device_controller/usbc_dsclen_6_s9  (
    .F(u_usb_device_controller_usbc_dsclen_6_14),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]),
    .I1(u_usb_device_controller_usbc_dsclen_6_16) 
);
defparam \u_usb_device_controller/usbc_dsclen_6_s9 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usbc_dsclen_6_s10  (
    .F(u_usb_device_controller_usbc_dsclen_6_15),
    .I0(desc_qual_len_i_d[6]),
    .I1(u_usb_device_controller_usbc_dsclen_6_17),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_6_s10 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/usbc_dsclen_7_s9  (
    .F(u_usb_device_controller_usbc_dsclen_7_14),
    .I0(u_usb_device_controller_usbc_dsclen_7_15),
    .I1(u_usb_device_controller_usbc_dsclen_7_16),
    .I2(u_usb_device_controller_usbc_dsclen_7_17),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_7_s9 .INIT=16'h0FBB;
  LUT4 \u_usb_device_controller/descrom_start_0_s9  (
    .F(u_usb_device_controller_descrom_start_0_14),
    .I0(desc_dev_addr_i_d[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_0_16),
    .I3(u_usb_device_controller_descrom_start_0_17) 
);
defparam \u_usb_device_controller/descrom_start_0_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_0_s10  (
    .F(u_usb_device_controller_descrom_start_0_15),
    .I0(u_usb_device_controller_descrom_start_0_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[0]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_0_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_1_s9  (
    .F(u_usb_device_controller_descrom_start_1_14),
    .I0(desc_dev_addr_i_d[1]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_1_16),
    .I3(u_usb_device_controller_descrom_start_1_17) 
);
defparam \u_usb_device_controller/descrom_start_1_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_1_s10  (
    .F(u_usb_device_controller_descrom_start_1_15),
    .I0(u_usb_device_controller_descrom_start_1_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[1]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_1_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_2_s9  (
    .F(u_usb_device_controller_descrom_start_2_14),
    .I0(desc_dev_addr_i_d[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_2_16),
    .I3(u_usb_device_controller_descrom_start_2_17) 
);
defparam \u_usb_device_controller/descrom_start_2_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_2_s10  (
    .F(u_usb_device_controller_descrom_start_2_15),
    .I0(u_usb_device_controller_descrom_start_2_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[2]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_2_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_3_s9  (
    .F(u_usb_device_controller_descrom_start_3_14),
    .I0(desc_dev_addr_i_d[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_3_16),
    .I3(u_usb_device_controller_descrom_start_3_17) 
);
defparam \u_usb_device_controller/descrom_start_3_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_3_s10  (
    .F(u_usb_device_controller_descrom_start_3_15),
    .I0(u_usb_device_controller_descrom_start_3_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[3]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_3_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_4_s9  (
    .F(u_usb_device_controller_descrom_start_4_14),
    .I0(desc_dev_addr_i_d[4]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_4_16),
    .I3(u_usb_device_controller_descrom_start_4_17) 
);
defparam \u_usb_device_controller/descrom_start_4_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_4_s10  (
    .F(u_usb_device_controller_descrom_start_4_15),
    .I0(u_usb_device_controller_descrom_start_4_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[4]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_4_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_5_s9  (
    .F(u_usb_device_controller_descrom_start_5_14),
    .I0(desc_dev_addr_i_d[5]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_5_16),
    .I3(u_usb_device_controller_descrom_start_5_17) 
);
defparam \u_usb_device_controller/descrom_start_5_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_5_s10  (
    .F(u_usb_device_controller_descrom_start_5_15),
    .I0(u_usb_device_controller_descrom_start_5_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[5]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_5_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_6_s9  (
    .F(u_usb_device_controller_descrom_start_6_14),
    .I0(desc_dev_addr_i_d[6]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_6_16),
    .I3(u_usb_device_controller_descrom_start_6_17) 
);
defparam \u_usb_device_controller/descrom_start_6_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_6_s10  (
    .F(u_usb_device_controller_descrom_start_6_15),
    .I0(u_usb_device_controller_descrom_start_6_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[6]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_6_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_7_s9  (
    .F(u_usb_device_controller_descrom_start_7_14),
    .I0(desc_dev_addr_i_d[7]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_7_16),
    .I3(u_usb_device_controller_descrom_start_7_17) 
);
defparam \u_usb_device_controller/descrom_start_7_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_7_s10  (
    .F(u_usb_device_controller_descrom_start_7_15),
    .I0(u_usb_device_controller_descrom_start_7_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[7]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_7_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_8_s9  (
    .F(u_usb_device_controller_descrom_start_8_14),
    .I0(desc_dev_addr_i_d[8]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_8_16),
    .I3(u_usb_device_controller_descrom_start_8_17) 
);
defparam \u_usb_device_controller/descrom_start_8_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_8_s10  (
    .F(u_usb_device_controller_descrom_start_8_15),
    .I0(u_usb_device_controller_descrom_start_8_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[8]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_8_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_9_s9  (
    .F(u_usb_device_controller_descrom_start_9_14),
    .I0(desc_dev_addr_i_d[9]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_descrom_start_9_16),
    .I3(u_usb_device_controller_descrom_start_9_17) 
);
defparam \u_usb_device_controller/descrom_start_9_s9 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/descrom_start_9_s10  (
    .F(u_usb_device_controller_descrom_start_9_15),
    .I0(u_usb_device_controller_descrom_start_9_18),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_addr_i_d[9]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/descrom_start_9_s10 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/usb_transact_inst/txpop_o_d_s1  (
    .F(u_usb_device_controller_usb_transact_inst_txpop_o_d_5),
    .I0(u_usb_device_controller_usb_transact_inst_n1157_27),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_28),
    .I2(u_usb_device_controller_usb_transact_inst_n1041_4),
    .I3(u_usb_device_controller_usb_transact_inst_txpop_o_d_7) 
);
defparam \u_usb_device_controller/usb_transact_inst/txpop_o_d_s1 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/test_packet_inst/n313_s4  (
    .F(u_usb_device_controller_test_packet_inst_n313_8),
    .I0(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I1(u_usb_device_controller_test_packet_inst_n313_9),
    .I2(u_usb_device_controller_test_packet_inst_cnt[5]),
    .I3(u_usb_device_controller_test_packet_inst_n318_9) 
);
defparam \u_usb_device_controller/test_packet_inst/n313_s4 .INIT=16'h1F00;
  LUT4 \u_usb_device_controller/test_packet_inst/n316_s4  (
    .F(u_usb_device_controller_test_packet_inst_n316_8),
    .I0(u_usb_device_controller_test_packet_inst_cnt[2]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I3(u_usb_device_controller_test_packet_inst_cnt_11_9) 
);
defparam \u_usb_device_controller/test_packet_inst/n316_s4 .INIT=16'hEF00;
  LUT3 \u_usb_device_controller/test_packet_inst/n314_s4  (
    .F(u_usb_device_controller_test_packet_inst_n314_8),
    .I0(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[2]) 
);
defparam \u_usb_device_controller/test_packet_inst/n314_s4 .INIT=8'h01;
  LUT4 \u_usb_device_controller/test_packet_inst/n314_s5  (
    .F(u_usb_device_controller_test_packet_inst_n314_9),
    .I0(u_usb_device_controller_test_packet_inst_n314_8),
    .I1(u_usb_device_controller_test_packet_inst_n133_7),
    .I2(u_usb_device_controller_test_packet_inst_n312_13),
    .I3(u_usb_device_controller_test_packet_inst_test_en_dly_Z) 
);
defparam \u_usb_device_controller/test_packet_inst/n314_s5 .INIT=16'h4F00;
  LUT2 \u_usb_device_controller/n1810_s2  (
    .F(u_usb_device_controller_n1810_6),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_s_osync) 
);
defparam \u_usb_device_controller/n1810_s2 .INIT=4'h6;
  LUT4 \u_usb_device_controller/u_usb_packet/n776_s2  (
    .F(u_usb_device_controller_u_usb_packet_n776_6),
    .I0(u_usb_device_controller_u_usb_packet_n774_7),
    .I1(u_usb_device_controller_u_usb_packet_n771_6),
    .I2(u_usb_device_controller_u_usb_packet_n770_6),
    .I3(u_usb_device_controller_u_usb_packet_n771_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n776_s2 .INIT=16'h6996;
  LUT2 \u_usb_device_controller/u_usb_packet/n776_s3  (
    .F(u_usb_device_controller_u_usb_packet_n776_7),
    .I0(u_usb_device_controller_u_usb_packet_n912_9),
    .I1(u_usb_device_controller_u_usb_packet_n767_6) 
);
defparam \u_usb_device_controller/u_usb_packet/n776_s3 .INIT=4'h6;
  LUT2 \u_usb_device_controller/u_usb_packet/n776_s4  (
    .F(u_usb_device_controller_u_usb_packet_n776_8),
    .I0(u_usb_device_controller_u_usb_packet_n774_6),
    .I1(u_usb_device_controller_u_usb_packet_n912_10) 
);
defparam \u_usb_device_controller/u_usb_packet/n776_s4 .INIT=4'h6;
  LUT2 \u_usb_device_controller/u_usb_packet/n776_s5  (
    .F(u_usb_device_controller_u_usb_packet_n776_9),
    .I0(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I1(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n776_s5 .INIT=4'h1;
  LUT2 \u_usb_device_controller/u_usb_packet/n775_s2  (
    .F(u_usb_device_controller_u_usb_packet_n775_6),
    .I0(u_usb_device_controller_u_usb_packet_n912_10),
    .I1(u_usb_device_controller_u_usb_packet_n771_6) 
);
defparam \u_usb_device_controller/u_usb_packet/n775_s2 .INIT=4'h6;
  LUT2 \u_usb_device_controller/u_usb_packet/n775_s3  (
    .F(u_usb_device_controller_u_usb_packet_n775_7),
    .I0(u_usb_device_controller_u_usb_packet_n912_9),
    .I1(u_usb_device_controller_u_usb_packet_n770_6) 
);
defparam \u_usb_device_controller/u_usb_packet/n775_s3 .INIT=4'h6;
  LUT3 \u_usb_device_controller/u_usb_packet/n775_s4  (
    .F(u_usb_device_controller_u_usb_packet_n775_8),
    .I0(u_usb_device_controller_u_usb_packet_n774_6),
    .I1(u_usb_device_controller_u_usb_packet_n767_6),
    .I2(u_usb_device_controller_u_usb_packet_n771_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n775_s4 .INIT=8'h96;
  LUT4 \u_usb_device_controller/u_usb_packet/n774_s2  (
    .F(u_usb_device_controller_u_usb_packet_n774_6),
    .I0(u_usb_device_controller_u_usb_packet_n642_21),
    .I1(u_usb_device_controller_u_usb_packet_n774_8),
    .I2(u_usb_device_controller_u_usb_packet_n774_9),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf[9]) 
);
defparam \u_usb_device_controller/u_usb_packet/n774_s2 .INIT=16'hF40B;
  LUT4 \u_usb_device_controller/u_usb_packet/n774_s3  (
    .F(u_usb_device_controller_u_usb_packet_n774_7),
    .I0(u_usb_device_controller_u_usb_packet_n640_21),
    .I1(u_usb_device_controller_u_usb_packet_n774_10),
    .I2(u_usb_device_controller_u_usb_packet_n774_11),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf[8]) 
);
defparam \u_usb_device_controller/u_usb_packet/n774_s3 .INIT=16'hF40B;
  LUT4 \u_usb_device_controller/u_usb_packet/n771_s2  (
    .F(u_usb_device_controller_u_usb_packet_n771_6),
    .I0(u_usb_device_controller_u_usb_packet_n646_20),
    .I1(u_usb_device_controller_u_usb_packet_n771_8),
    .I2(u_usb_device_controller_u_usb_packet_n771_9),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf[11]) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s2 .INIT=16'hF40B;
  LUT4 \u_usb_device_controller/u_usb_packet/n771_s3  (
    .F(u_usb_device_controller_u_usb_packet_n771_7),
    .I0(u_usb_device_controller_u_usb_packet_n771_10),
    .I1(u_usb_device_controller_u_usb_packet_n771_11),
    .I2(u_usb_device_controller_u_usb_packet_n771_12),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf[12]) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s3 .INIT=16'hF40B;
  LUT4 \u_usb_device_controller/u_usb_packet/n770_s2  (
    .F(u_usb_device_controller_u_usb_packet_n770_6),
    .I0(u_usb_device_controller_u_usb_packet_n650_20),
    .I1(u_usb_device_controller_u_usb_packet_n770_12),
    .I2(u_usb_device_controller_u_usb_packet_n770_10),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf[13]) 
);
defparam \u_usb_device_controller/u_usb_packet/n770_s2 .INIT=16'hF40B;
  LUT4 \u_usb_device_controller/u_usb_packet/n767_s2  (
    .F(u_usb_device_controller_u_usb_packet_n767_6),
    .I0(u_usb_device_controller_u_usb_packet_n328_16),
    .I1(u_usb_device_controller_u_usb_packet_n767_12),
    .I2(u_usb_device_controller_u_usb_packet_n767_8),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf[15]) 
);
defparam \u_usb_device_controller/u_usb_packet/n767_s2 .INIT=16'h8F70;
  LUT3 \u_usb_device_controller/u_usb_packet/n761_s2  (
    .F(u_usb_device_controller_u_usb_packet_n761_6),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[7]),
    .I1(u_usb_device_controller_u_usb_packet_n767_6),
    .I2(u_usb_device_controller_u_usb_packet_n912_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n761_s2 .INIT=8'h96;
  LUT4 \u_usb_device_controller/u_usb_init/n217_s28  (
    .F(u_usb_device_controller_u_usb_init_n217_37),
    .I0(u_usb_device_controller_u_usb_init_s_state[2]),
    .I1(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_u_usb_init_s_linestate[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n217_s28 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/u_usb_init/n217_s29  (
    .F(u_usb_device_controller_u_usb_init_n217_38),
    .I0(u_usb_device_controller_u_usb_init_s_state[1]),
    .I1(u_usb_device_controller_u_usb_init_s_state[2]) 
);
defparam \u_usb_device_controller/u_usb_init/n217_s29 .INIT=4'h1;
  LUT4 \u_usb_device_controller/usb_control_inst/usbc_dscrd_s0  (
    .F(u_usb_device_controller_usb_control_inst_usbc_dscrd_4),
    .I0(u_usb_device_controller_usb_control_inst_s_state[8]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1661_22) 
);
defparam \u_usb_device_controller/usb_control_inst/usbc_dscrd_s0 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/s_answerptr_7_s9  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_7_13),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I1(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[9]),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_7_11) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_7_s9 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s10  (
    .F(u_usb_device_controller_usb_control_inst_s_sendbyte_7_14),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s10 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_control_inst/s_interface_set_s5  (
    .F(u_usb_device_controller_usb_control_inst_s_interface_set_8),
    .I0(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_11) 
);
defparam \u_usb_device_controller/usb_control_inst/s_interface_set_s5 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_control_inst/s_interface_set_s6  (
    .F(u_usb_device_controller_usb_control_inst_s_interface_set_9),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I1(u_usb_device_controller_usb_control_inst_n1837_6),
    .I2(u_usb_device_controller_usb_control_inst_n1876_13) 
);
defparam \u_usb_device_controller/usb_control_inst/s_interface_set_s6 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1133_s20  (
    .F(u_usb_device_controller_usb_transact_inst_n1133_26),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[9]),
    .I1(u_usb_device_controller_usb_transact_inst_n1146_22),
    .I2(u_usb_device_controller_usb_transact_inst_n1133_27),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_31) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1133_s20 .INIT=16'h4000;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1127_s20  (
    .F(u_usb_device_controller_usb_transact_inst_n1127_26),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[10]),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[11]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1127_s20 .INIT=4'h1;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1118_s20  (
    .F(u_usb_device_controller_usb_transact_inst_n1118_26),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[13]),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[14]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1118_s20 .INIT=4'h1;
  LUT2 \u_usb_device_controller/n1613_s15  (
    .F(u_usb_device_controller_n1613_21),
    .I0(u_usb_device_controller_n1585),
    .I1(u_usb_device_controller_n1615_15) 
);
defparam \u_usb_device_controller/n1613_s15 .INIT=4'h1;
  LUT2 \u_usb_device_controller/n1611_s15  (
    .F(u_usb_device_controller_n1611_21),
    .I0(u_usb_device_controller_s_bufptr[0]),
    .I1(u_usb_device_controller_s_bufptr[1]) 
);
defparam \u_usb_device_controller/n1611_s15 .INIT=4'h8;
  LUT2 \u_usb_device_controller/n1603_s15  (
    .F(u_usb_device_controller_n1603_21),
    .I0(u_usb_device_controller_s_bufptr[4]),
    .I1(u_usb_device_controller_s_bufptr[5]) 
);
defparam \u_usb_device_controller/n1603_s15 .INIT=4'h8;
  LUT2 \u_usb_device_controller/n1597_s15  (
    .F(u_usb_device_controller_n1597_21),
    .I0(u_usb_device_controller_s_bufptr[7]),
    .I1(u_usb_device_controller_s_bufptr[8]) 
);
defparam \u_usb_device_controller/n1597_s15 .INIT=4'h8;
  LUT4 \u_usb_device_controller/u_usb_packet/n579_s13  (
    .F(u_usb_device_controller_u_usb_packet_n579_19),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf[3]),
    .I2(u_usb_device_controller_u_usb_packet_n579_21),
    .I3(u_usb_device_controller_u_usb_packet_n579_22) 
);
defparam \u_usb_device_controller/u_usb_packet/n579_s13 .INIT=16'h6996;
  LUT4 \u_usb_device_controller/u_usb_packet/n579_s14  (
    .F(u_usb_device_controller_u_usb_packet_n579_20),
    .I0(u_usb_device_controller_u_usb_packet_s_state[3]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[2]),
    .I2(u_usb_device_controller_u_usb_packet_n784_9),
    .I3(u_usb_device_controller_u_usb_packet_n784_11) 
);
defparam \u_usb_device_controller/u_usb_packet/n579_s14 .INIT=16'h4000;
  LUT3 \u_usb_device_controller/u_usb_packet/n577_s13  (
    .F(u_usb_device_controller_u_usb_packet_n577_19),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf[1]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]) 
);
defparam \u_usb_device_controller/u_usb_packet/n577_s13 .INIT=8'h96;
  LUT4 \u_usb_device_controller/u_usb_packet/n577_s14  (
    .F(u_usb_device_controller_u_usb_packet_n577_20),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf[4]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I3(u_usb_device_controller_u_usb_packet_crc5_buf[3]) 
);
defparam \u_usb_device_controller/u_usb_packet/n577_s14 .INIT=16'h6996;
  LUT4 \u_usb_device_controller/u_usb_packet/n575_s13  (
    .F(u_usb_device_controller_u_usb_packet_n575_19),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf[0]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]) 
);
defparam \u_usb_device_controller/u_usb_packet/n575_s13 .INIT=16'h6996;
  LUT4 \u_usb_device_controller/u_usb_packet/n573_s13  (
    .F(u_usb_device_controller_u_usb_packet_n573_19),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf[4]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .I3(u_usb_device_controller_u_usb_packet_crc5_buf[0]) 
);
defparam \u_usb_device_controller/u_usb_packet/n573_s13 .INIT=16'h6996;
  LUT4 \u_usb_device_controller/u_usb_packet/n571_s13  (
    .F(u_usb_device_controller_u_usb_packet_n571_19),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf[1]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I3(u_usb_device_controller_u_usb_packet_n579_21) 
);
defparam \u_usb_device_controller/u_usb_packet/n571_s13 .INIT=16'h6996;
  LUT3 \u_usb_device_controller/utmi_dataout_o_d_7_s3  (
    .F(u_usb_device_controller_utmi_dataout_o_d_7_7),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_utmi_dataout_o_d_0_4) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_7_s3 .INIT=8'h40;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_0_s1  (
    .F(u_usb_device_controller_utmi_dataout_o_d_0_4),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[6]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_testmode[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_testmode[1]),
    .I3(u_usb_device_controller_utmi_dataout_o_d_7_8) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_0_s1 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/utmi_dataout_o_d_0_s2  (
    .F(u_usb_device_controller_utmi_dataout_o_d_0_5),
    .I0(u_usb_device_controller_test_packet_inst_test_data_Z[0]),
    .I1(u_usb_device_controller_u_usb_packet_usbp_dataout_o[0]),
    .I2(u_usb_device_controller_test_packet_inst_cnt_11_10) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_0_s2 .INIT=8'hAC;
  LUT4 \u_usb_device_controller/n2339_s2  (
    .F(u_usb_device_controller_n2339_5),
    .I0(txdat_len_i_d[6]),
    .I1(txdat_len_i_d[7]),
    .I2(txdat_len_i_d[8]),
    .I3(txdat_len_i_d[9]) 
);
defparam \u_usb_device_controller/n2339_s2 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/n2339_s3  (
    .F(u_usb_device_controller_n2339_6),
    .I0(txdat_len_i_d[2]),
    .I1(txdat_len_i_d[3]),
    .I2(txdat_len_i_d[4]),
    .I3(txdat_len_i_d[5]) 
);
defparam \u_usb_device_controller/n2339_s3 .INIT=16'h0001;
  LUT2 \u_usb_device_controller/n2024_s2  (
    .F(u_usb_device_controller_n2024_5),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]),
    .I1(u_usb_device_controller_n2024_7) 
);
defparam \u_usb_device_controller/n2024_s2 .INIT=4'h4;
  LUT4 \u_usb_device_controller/n2024_s3  (
    .F(u_usb_device_controller_n2024_6),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[7]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/n2024_s3 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/test_packet_inst/n130_s4  (
    .F(u_usb_device_controller_test_packet_inst_n130_7),
    .I0(u_usb_device_controller_test_packet_inst_cnt[6]),
    .I1(u_usb_device_controller_test_packet_inst_cnt_11_11),
    .I2(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I3(u_usb_device_controller_test_packet_inst_n318_13) 
);
defparam \u_usb_device_controller/test_packet_inst/n130_s4 .INIT=16'h7F00;
  LUT4 \u_usb_device_controller/test_packet_inst/n378_s2  (
    .F(u_usb_device_controller_test_packet_inst_n378_5),
    .I0(u_usb_device_controller_test_packet_inst_cnt[6]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[7]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[8]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[9]) 
);
defparam \u_usb_device_controller/test_packet_inst/n378_s2 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/u_usb_packet/n782_s3  (
    .F(u_usb_device_controller_u_usb_packet_n782_6),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[3]),
    .I2(u_usb_device_controller_u_usb_packet_n640_27),
    .I3(u_usb_device_controller_u_usb_packet_n771_10) 
);
defparam \u_usb_device_controller/u_usb_packet/n782_s3 .INIT=16'h000E;
  LUT4 \u_usb_device_controller/u_usb_packet/n782_s4  (
    .F(u_usb_device_controller_u_usb_packet_n782_7),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[4]),
    .I1(u_usb_device_controller_u_usb_packet_n620),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf[12]),
    .I3(u_usb_device_controller_u_usb_packet_n622) 
);
defparam \u_usb_device_controller/u_usb_packet/n782_s4 .INIT=16'hB0BB;
  LUT4 \u_usb_device_controller/u_usb_packet/n782_s5  (
    .F(u_usb_device_controller_u_usb_packet_n782_8),
    .I0(u_usb_device_controller_u_usb_packet_s_txfirst),
    .I1(u_usb_device_controller_u_usb_packet_n615_49),
    .I2(u_usb_device_controller_u_usb_packet_n620_47),
    .I3(u_usb_device_controller_u_usb_packet_s_txready) 
);
defparam \u_usb_device_controller/u_usb_packet/n782_s5 .INIT=16'h00F4;
  LUT4 \u_usb_device_controller/u_usb_packet/n782_s6  (
    .F(u_usb_device_controller_u_usb_packet_n782_9),
    .I0(u_usb_device_controller_u_usb_packet_n626_42),
    .I1(u_usb_device_controller_u_usb_packet_n919_5),
    .I2(u_usb_device_controller_u_usb_packet_n626_46),
    .I3(u_usb_device_controller_u_usb_packet_n784_18) 
);
defparam \u_usb_device_controller/u_usb_packet/n782_s6 .INIT=16'h4F00;
  LUT4 \u_usb_device_controller/u_usb_packet/n784_s4  (
    .F(u_usb_device_controller_u_usb_packet_n784_7),
    .I0(u_usb_device_controller_u_usb_packet_n328_12),
    .I1(u_usb_device_controller_u_usb_packet_n328_13),
    .I2(u_usb_device_controller_u_usb_packet_n328_14),
    .I3(u_usb_device_controller_u_usb_packet_n784_13) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s4 .INIT=16'h4F00;
  LUT4 \u_usb_device_controller/u_usb_packet/n784_s5  (
    .F(u_usb_device_controller_u_usb_packet_n784_8),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[6]),
    .I1(u_usb_device_controller_u_usb_packet_n620),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout[1]),
    .I3(u_usb_device_controller_u_usb_packet_n782_8) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s5 .INIT=16'h0BBB;
  LUT3 \u_usb_device_controller/u_usb_packet/n784_s6  (
    .F(u_usb_device_controller_u_usb_packet_n784_9),
    .I0(u_usb_device_controller_u_usb_packet_s_state[4]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[5]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[6]) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s6 .INIT=8'h01;
  LUT2 \u_usb_device_controller/u_usb_packet/n784_s7  (
    .F(u_usb_device_controller_u_usb_packet_n784_10),
    .I0(u_usb_device_controller_u_usb_packet_s_state[2]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[3]) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s7 .INIT=4'h1;
  LUT4 \u_usb_device_controller/u_usb_packet/n784_s8  (
    .F(u_usb_device_controller_u_usb_packet_n784_11),
    .I0(u_usb_device_controller_u_usb_packet_s_state[0]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[1]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[7]),
    .I3(u_usb_device_controller_u_usb_packet_s_state[8]) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s8 .INIT=16'h0001;
  LUT3 \u_usb_device_controller/u_usb_packet/n785_s3  (
    .F(u_usb_device_controller_u_usb_packet_n785_6),
    .I0(u_usb_device_controller_u_usb_packet_n919_5),
    .I1(u_usb_device_controller_u_usb_packet_n626_42),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54) 
);
defparam \u_usb_device_controller/u_usb_packet/n785_s3 .INIT=8'hD0;
  LUT3 \u_usb_device_controller/u_usb_packet/n785_s4  (
    .F(u_usb_device_controller_u_usb_packet_n785_7),
    .I0(u_usb_device_controller_u_usb_packet_n622),
    .I1(u_usb_device_controller_u_usb_packet_crc16_buf[15]),
    .I2(u_usb_device_controller_u_usb_packet_n785_8) 
);
defparam \u_usb_device_controller/u_usb_packet/n785_s4 .INIT=8'hD0;
  LUT4 \u_usb_device_controller/u_usb_packet/n1454_s2  (
    .F(u_usb_device_controller_u_usb_packet_n1454_5),
    .I0(u_usb_device_controller_u_usb_packet_s_state[7]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[8]),
    .I2(u_usb_device_controller_u_usb_packet_n784_9),
    .I3(u_usb_device_controller_u_usb_packet_n784_10) 
);
defparam \u_usb_device_controller/u_usb_packet/n1454_s2 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/u_usb_packet/n912_s5  (
    .F(u_usb_device_controller_u_usb_packet_n912_8),
    .I0(u_usb_device_controller_u_usb_packet_n912_14),
    .I1(u_usb_device_controller_u_usb_packet_n912_15) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s5 .INIT=4'h8;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s6  (
    .F(u_usb_device_controller_u_usb_packet_n912_9),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I1(u_usb_device_controller_u_usb_packet_n785_6),
    .I2(u_usb_device_controller_u_usb_packet_n784_7),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf[14]) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s6 .INIT=16'hF20D;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s7  (
    .F(u_usb_device_controller_u_usb_packet_n912_10),
    .I0(u_usb_device_controller_u_usb_packet_n644_21),
    .I1(u_usb_device_controller_u_usb_packet_n912_16),
    .I2(u_usb_device_controller_u_usb_packet_n912_17),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf[10]) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s7 .INIT=16'hF40B;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s8  (
    .F(u_usb_device_controller_u_usb_packet_n912_11),
    .I0(u_usb_device_controller_u_usb_packet_n912_18),
    .I1(u_usb_device_controller_u_usb_packet_n571_19),
    .I2(u_usb_device_controller_u_usb_packet_n912_19),
    .I3(u_usb_device_controller_u_usb_packet_n628) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s8 .INIT=16'h00EF;
  LUT3 \u_usb_device_controller/u_usb_packet/n912_s9  (
    .F(u_usb_device_controller_u_usb_packet_n912_12),
    .I0(u_usb_device_controller_u_usb_packet_n912_20),
    .I1(u_usb_device_controller_u_usb_packet_n912_21),
    .I2(u_usb_device_controller_u_usb_packet_s_rxgoodpacket) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s9 .INIT=8'hB0;
  LUT3 \u_usb_device_controller/u_usb_packet/n912_s10  (
    .F(u_usb_device_controller_u_usb_packet_n912_13),
    .I0(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I1(u_usb_device_controller_u_usb_packet_n785_6),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf_15_14) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s10 .INIT=8'h01;
  LUT3 \u_usb_device_controller/u_usb_packet/n919_s2  (
    .F(u_usb_device_controller_u_usb_packet_n919_5),
    .I0(u_usb_device_controller_usb_transact_inst_n1072_18),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[5]),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_50) 
);
defparam \u_usb_device_controller/u_usb_packet/n919_s2 .INIT=8'h07;
  LUT3 \u_usb_device_controller/u_usb_packet/n920_s3  (
    .F(u_usb_device_controller_u_usb_packet_n920_6),
    .I0(u_usb_device_controller_u_usb_packet_s_state[7]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[8]),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout_7_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n920_s3 .INIT=8'h40;
  LUT3 \u_usb_device_controller/u_usb_packet/n920_s4  (
    .F(u_usb_device_controller_u_usb_packet_n920_7),
    .I0(u_usb_device_controller_u_usb_packet_n615_49),
    .I1(u_usb_device_controller_u_usb_packet_n620_47),
    .I2(u_usb_device_controller_u_usb_packet_n800_6) 
);
defparam \u_usb_device_controller/u_usb_packet/n920_s4 .INIT=8'h01;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1565_s4  (
    .F(u_usb_device_controller_usb_transact_inst_n1565_7),
    .I0(u_usb_device_controller_usb_transact_inst_s_out),
    .I1(u_usb_device_controller_usb_transact_inst_s_setup_2),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1565_s4 .INIT=16'h0E00;
  LUT4 \u_usb_device_controller/usb_control_inst/n2902_s2  (
    .F(u_usb_device_controller_usb_control_inst_n2902_5),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I3(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n2902_s2 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/u_usb_init/n212_s25  (
    .F(u_usb_device_controller_u_usb_init_n212_33),
    .I0(u_usb_device_controller_u_usb_init_s_state_3_12),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s25 .INIT=4'h4;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s27  (
    .F(u_usb_device_controller_u_usb_init_n212_35),
    .I0(u_usb_device_controller_u_usb_init_s_chirpcnt[1]),
    .I1(u_usb_device_controller_u_usb_init_s_chirpcnt[0]),
    .I2(u_usb_device_controller_u_usb_init_s_chirpcnt[2]),
    .I3(u_usb_device_controller_u_usb_init_s_chirpcnt_2_9) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s27 .INIT=16'h4000;
  LUT3 \u_usb_device_controller/u_usb_init/n212_s29  (
    .F(u_usb_device_controller_u_usb_init_n212_37),
    .I0(u_usb_device_controller_u_usb_init_n216_53),
    .I1(u_usb_device_controller_u_usb_init_s_chirpcnt_2_10),
    .I2(u_usb_device_controller_u_usb_init_n212_44) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s29 .INIT=8'h01;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s30  (
    .F(u_usb_device_controller_u_usb_init_n212_38),
    .I0(u_usb_device_controller_u_usb_init_s_linestate[1]),
    .I1(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .I2(u_usb_device_controller_u_usb_init_n212_45),
    .I3(u_usb_device_controller_u_usb_init_s_state[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s30 .INIT=16'hBBF0;
  LUT2 \u_usb_device_controller/u_usb_init/n212_s31  (
    .F(u_usb_device_controller_u_usb_init_n212_39),
    .I0(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I1(u_usb_device_controller_u_usb_init_s_state[3]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s31 .INIT=4'h1;
  LUT2 \u_usb_device_controller/u_usb_init/n215_s46  (
    .F(u_usb_device_controller_u_usb_init_n215_53),
    .I0(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .I1(u_usb_device_controller_u_usb_init_s_linestate[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s46 .INIT=4'h1;
  LUT3 \u_usb_device_controller/u_usb_init/n215_s47  (
    .F(u_usb_device_controller_u_usb_init_n215_54),
    .I0(u_usb_device_controller_u_usb_init_n215_58),
    .I1(u_usb_device_controller_u_usb_init_n215_59),
    .I2(u_usb_device_controller_u_usb_init_n215_67) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s47 .INIT=8'h80;
  LUT4 \u_usb_device_controller/u_usb_init/n215_s50  (
    .F(u_usb_device_controller_u_usb_init_n215_57),
    .I0(u_usb_device_controller_u_usb_init_s_state[1]),
    .I1(u_usb_device_controller_u_usb_init_n212_44),
    .I2(u_usb_device_controller_u_usb_init_s_state[2]),
    .I3(u_usb_device_controller_u_usb_init_s_state[3]) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s50 .INIT=16'h00EF;
  LUT2 \u_usb_device_controller/u_usb_init/n216_s46  (
    .F(u_usb_device_controller_u_usb_init_n216_52),
    .I0(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4) 
);
defparam \u_usb_device_controller/u_usb_init/n216_s46 .INIT=4'h8;
  LUT3 \u_usb_device_controller/u_usb_init/n216_s47  (
    .F(u_usb_device_controller_u_usb_init_n216_53),
    .I0(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I1(u_usb_device_controller_u_usb_init_n212_41),
    .I2(u_usb_device_controller_u_usb_init_n212_42) 
);
defparam \u_usb_device_controller/u_usb_init/n216_s47 .INIT=8'h40;
  LUT3 \u_usb_device_controller/u_usb_init/n216_s48  (
    .F(u_usb_device_controller_u_usb_init_n216_54),
    .I0(u_usb_device_controller_u_usb_init_s_chirpcnt_2_10),
    .I1(u_usb_device_controller_u_usb_init_s_state[3]),
    .I2(u_usb_device_controller_u_usb_init_n215_57) 
);
defparam \u_usb_device_controller/u_usb_init/n216_s48 .INIT=8'h0D;
  LUT3 \u_usb_device_controller/usb_control_inst/n435_s14  (
    .F(u_usb_device_controller_usb_control_inst_n435_18),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_n1864_8) 
);
defparam \u_usb_device_controller/usb_control_inst/n435_s14 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n435_s15  (
    .F(u_usb_device_controller_usb_control_inst_n435_19),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I3(u_usb_device_controller_usb_control_inst_n1836_10) 
);
defparam \u_usb_device_controller/usb_control_inst/n435_s15 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/usb_control_inst/n435_s16  (
    .F(u_usb_device_controller_usb_control_inst_n435_20),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n435_s16 .INIT=4'h1;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s8  (
    .F(u_usb_device_controller_u_usb_packet_n328_12),
    .I0(u_usb_device_controller_usb_transact_inst_n1080_46),
    .I1(u_usb_device_controller_usb_transact_inst_n1138_25),
    .I2(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_5_10) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s8 .INIT=16'h7000;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s9  (
    .F(u_usb_device_controller_u_usb_packet_n328_13),
    .I0(u_usb_device_controller_u_usb_packet_n328_20),
    .I1(descrom_rdata_i_d[1]),
    .I2(u_usb_device_controller_usb_control_inst_n1649_18),
    .I3(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s9 .INIT=16'hCA00;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s10  (
    .F(u_usb_device_controller_u_usb_packet_n328_14),
    .I0(u_usb_device_controller_usb_transact_inst_n1080_46),
    .I1(u_usb_device_controller_usb_transact_inst_n1138_25),
    .I2(u_usb_device_controller_u_usb_packet_n328_21),
    .I3(u_usb_device_controller_u_usb_packet_n328_22) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s10 .INIT=16'h8F00;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s12  (
    .F(u_usb_device_controller_u_usb_packet_n328_16),
    .I0(u_usb_device_controller_u_usb_packet_n328_23),
    .I1(descrom_rdata_i_d[0]),
    .I2(u_usb_device_controller_usb_control_inst_n1649_18),
    .I3(u_usb_device_controller_u_usb_packet_n328_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s12 .INIT=16'hCCCA;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s13  (
    .F(u_usb_device_controller_u_usb_packet_n328_17),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[0]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[1]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s13 .INIT=16'h0001;
  LUT2 \u_usb_device_controller/usb_control_inst/n1836_s6  (
    .F(u_usb_device_controller_usb_control_inst_n1836_9),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I1(u_usb_device_controller_usb_control_inst_n1836_11) 
);
defparam \u_usb_device_controller/usb_control_inst/n1836_s6 .INIT=4'h4;
  LUT3 \u_usb_device_controller/usb_control_inst/n1836_s7  (
    .F(u_usb_device_controller_usb_control_inst_n1836_10),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I1(u_usb_device_controller_usb_control_inst_n1836_11),
    .I2(u_usb_device_controller_usb_control_inst_n1715_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1836_s7 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_endpt_0_s4  (
    .F(u_usb_device_controller_usb_transact_inst_s_endpt_0_7),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[0]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[3]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[1]),
    .I3(u_usb_device_controller_usb_transact_inst_n1074_25) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_endpt_0_s4 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/u_usb_init/s_state_3_s6  (
    .F(u_usb_device_controller_u_usb_init_s_state_3_11),
    .I0(u_usb_device_controller_u_usb_init_s_state_3_12),
    .I1(u_usb_device_controller_u_usb_init_n212_57) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s6 .INIT=4'h1;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_3_s7  (
    .F(u_usb_device_controller_u_usb_init_s_state_3_12),
    .I0(u_usb_device_controller_u_usb_init_s_state_3_13),
    .I1(u_usb_device_controller_u_usb_init_n215_59),
    .I2(u_usb_device_controller_u_usb_init_s_state_3_14),
    .I3(u_usb_device_controller_u_usb_init_s_state_3_18) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s7 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s5  (
    .F(u_usb_device_controller_u_usb_init_s_chirpcnt_2_9),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[0]),
    .I1(u_usb_device_controller_u_usb_init_n212_41),
    .I2(u_usb_device_controller_u_usb_init_s_chirpcnt_2_11),
    .I3(u_usb_device_controller_u_usb_init_s_chirpcnt_2_12) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s5 .INIT=16'h8000;
  LUT3 \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s6  (
    .F(u_usb_device_controller_u_usb_init_s_chirpcnt_2_10),
    .I0(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I1(u_usb_device_controller_u_usb_init_s_chirpcnt_2_13),
    .I2(u_usb_device_controller_u_usb_init_s_chirpcnt_2_14) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s6 .INIT=8'h80;
  LUT3 \u_usb_device_controller/u_usb_packet/n615_s39  (
    .F(u_usb_device_controller_u_usb_packet_n615_43),
    .I0(u_usb_device_controller_u_usb_packet_s_state[4]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[5]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[6]) 
);
defparam \u_usb_device_controller/u_usb_packet/n615_s39 .INIT=8'h10;
  LUT4 \u_usb_device_controller/u_usb_packet/n615_s40  (
    .F(u_usb_device_controller_u_usb_packet_n615_44),
    .I0(u_usb_device_controller_u_usb_packet_s_state[5]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[6]),
    .I2(u_usb_device_controller_u_usb_packet_n615_47),
    .I3(u_usb_device_controller_u_usb_packet_n784_11) 
);
defparam \u_usb_device_controller/u_usb_packet/n615_s40 .INIT=16'h0100;
  LUT3 \u_usb_device_controller/u_usb_packet/n615_s41  (
    .F(u_usb_device_controller_u_usb_packet_n615_45),
    .I0(u_usb_device_controller_u_usb_packet_s_state[8]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[7]),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout_7_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n615_s41 .INIT=8'h70;
  LUT3 \u_usb_device_controller/u_usb_packet/n615_s42  (
    .F(u_usb_device_controller_u_usb_packet_n615_46),
    .I0(u_usb_device_controller_u_usb_packet_s_state[0]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[1]),
    .I2(u_usb_device_controller_u_usb_packet_n1454_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n615_s42 .INIT=8'h60;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1080_s44  (
    .F(u_usb_device_controller_usb_transact_inst_n1080_48),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[1]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[2]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[3]),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[0]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1080_s44 .INIT=16'h0100;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1080_s45  (
    .F(u_usb_device_controller_usb_transact_inst_n1080_49),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[11]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[12]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1080_s45 .INIT=8'hE9;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1064_s15  (
    .F(u_usb_device_controller_usb_transact_inst_n1064_20),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[11]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[12]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[10]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1064_s15 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1074_s20  (
    .F(u_usb_device_controller_usb_transact_inst_n1074_25),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[2]),
    .I1(u_usb_device_controller_usb_transact_inst_n1041_4),
    .I2(u_usb_device_controller_usb_transact_inst_n1041_8) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1074_s20 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1072_s15  (
    .F(u_usb_device_controller_usb_transact_inst_n1072_21),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[6]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[9]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1072_s15 .INIT=16'h0001;
  LUT3 \u_usb_device_controller/usb_control_inst/n1670_s39  (
    .F(u_usb_device_controller_usb_control_inst_n1670_43),
    .I0(u_usb_device_controller_usb_control_inst_s_state[1]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_15) 
);
defparam \u_usb_device_controller/usb_control_inst/n1670_s39 .INIT=8'h40;
  LUT3 \u_usb_device_controller/usb_control_inst/s_answerptr_7_s10  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_7_14),
    .I0(u_usb_device_controller_usb_control_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[5]),
    .I2(u_usb_device_controller_usb_control_inst_n1629_4) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_7_s10 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_control_inst/s_answerptr_7_s11  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_7_15),
    .I0(u_usb_device_controller_usb_control_inst_s_state[2]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[3]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_16) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_7_s11 .INIT=8'h10;
  LUT3 \u_usb_device_controller/usb_control_inst/s_answerptr_5_s9  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_5_12),
    .I0(u_usb_device_controller_usb_control_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[5]) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_5_s9 .INIT=8'h10;
  LUT4 \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s11  (
    .F(u_usb_device_controller_usb_control_inst_s_sendbyte_7_15),
    .I0(u_usb_device_controller_u_usb_packet_n800_6),
    .I1(u_usb_device_controller_u_usb_packet_n785_6),
    .I2(u_usb_device_controller_usb_transact_inst_txpop_o_d_5),
    .I3(u_usb_device_controller_usb_control_inst_n1672_44) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s11 .INIT=16'hE000;
  LUT4 \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s12  (
    .F(u_usb_device_controller_usb_control_inst_s_sendbyte_7_16),
    .I0(u_usb_device_controller_usb_control_inst_n1836_15),
    .I1(u_usb_device_controller_usb_control_inst_n1837_7),
    .I2(u_usb_device_controller_usb_control_inst_s_sendbyte_7_17),
    .I3(u_usb_device_controller_usb_control_inst_n1864_8) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s12 .INIT=16'hF800;
  LUT3 \u_usb_device_controller/u_usb_packet/s_state_11_s16  (
    .F(u_usb_device_controller_u_usb_packet_s_state_11_21),
    .I0(u_usb_device_controller_u_usb_packet_n784_20),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I2(u_usb_device_controller_u_usb_packet_s_state_11_27) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_11_s16 .INIT=8'h0D;
  LUT2 \u_usb_device_controller/u_usb_packet/s_state_11_s17  (
    .F(u_usb_device_controller_u_usb_packet_s_state_11_22),
    .I0(u_usb_device_controller_u_usb_init_usbp_chirpk),
    .I1(u_usb_device_controller_u_usb_packet_n784_18) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_11_s17 .INIT=4'h4;
  LUT4 \u_usb_device_controller/u_usb_packet/s_state_11_s18  (
    .F(u_usb_device_controller_u_usb_packet_s_state_11_23),
    .I0(u_usb_device_controller_u_usb_packet_n920_9),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf_4_13),
    .I2(u_usb_device_controller_u_usb_packet_n912_21),
    .I3(u_usb_device_controller_u_usb_packet_s_state_11_25) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_11_s18 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s8  (
    .F(u_usb_device_controller_usb_transact_inst_s_sendpid_3_13),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid_3_16) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s8 .INIT=4'h4;
  LUT3 \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s9  (
    .F(u_usb_device_controller_usb_transact_inst_s_sendpid_3_14),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3_17),
    .I1(u_usb_device_controller_usb_control_inst_n1670_43),
    .I2(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s9 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/u_usb_packet/n640_s16  (
    .F(u_usb_device_controller_u_usb_packet_n640_21),
    .I0(u_usb_device_controller_u_usb_packet_n328_12),
    .I1(u_usb_device_controller_usb_control_inst_n1649_18),
    .I2(u_usb_device_controller_u_usb_packet_n640_22),
    .I3(u_usb_device_controller_u_usb_packet_n640_23) 
);
defparam \u_usb_device_controller/u_usb_packet/n640_s16 .INIT=16'hEF00;
  LUT4 \u_usb_device_controller/u_usb_packet/n642_s16  (
    .F(u_usb_device_controller_u_usb_packet_n642_21),
    .I0(u_usb_device_controller_u_usb_packet_n328_12),
    .I1(u_usb_device_controller_usb_control_inst_n1649_18),
    .I2(u_usb_device_controller_u_usb_packet_n642_22),
    .I3(u_usb_device_controller_u_usb_packet_n642_23) 
);
defparam \u_usb_device_controller/u_usb_packet/n642_s16 .INIT=16'hEF00;
  LUT3 \u_usb_device_controller/u_usb_packet/n644_s16  (
    .F(u_usb_device_controller_u_usb_packet_n644_21),
    .I0(u_usb_device_controller_u_usb_packet_n644_22),
    .I1(u_usb_device_controller_u_usb_packet_n328_12),
    .I2(u_usb_device_controller_u_usb_packet_n644_23) 
);
defparam \u_usb_device_controller/u_usb_packet/n644_s16 .INIT=8'hD0;
  LUT4 \u_usb_device_controller/u_usb_packet/n646_s15  (
    .F(u_usb_device_controller_u_usb_packet_n646_20),
    .I0(u_usb_device_controller_u_usb_packet_n646_21),
    .I1(u_usb_device_controller_u_usb_packet_n328_12),
    .I2(u_usb_device_controller_u_usb_packet_n646_22),
    .I3(u_usb_device_controller_u_usb_packet_n646_23) 
);
defparam \u_usb_device_controller/u_usb_packet/n646_s15 .INIT=16'h10D0;
  LUT3 \u_usb_device_controller/u_usb_packet/n650_s15  (
    .F(u_usb_device_controller_u_usb_packet_n650_20),
    .I0(u_usb_device_controller_u_usb_packet_n328_12),
    .I1(u_usb_device_controller_u_usb_packet_n650_22),
    .I2(u_usb_device_controller_u_usb_packet_n650_23) 
);
defparam \u_usb_device_controller/u_usb_packet/n650_s15 .INIT=8'h10;
  LUT4 \u_usb_device_controller/u_usb_packet/n650_s16  (
    .F(u_usb_device_controller_u_usb_packet_n650_21),
    .I0(u_usb_device_controller_u_usb_packet_n650_23),
    .I1(u_usb_device_controller_u_usb_packet_n650_24),
    .I2(u_usb_device_controller_usb_transact_inst_s_sendpid[2]),
    .I3(u_usb_device_controller_u_usb_packet_n919_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n650_s16 .INIT=16'h7770;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1064_s16  (
    .F(u_usb_device_controller_usb_transact_inst_n1064_21),
    .I0(u_usb_device_controller_usb_transact_inst_n1068_18),
    .I1(u_usb_device_controller_usb_transact_inst_n1088_48) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1064_s16 .INIT=4'h8;
  LUT3 \u_usb_device_controller/usb_control_inst/n1672_s41  (
    .F(u_usb_device_controller_usb_control_inst_n1672_45),
    .I0(u_usb_device_controller_usb_control_inst_n1672_47),
    .I1(u_usb_device_controller_usb_control_inst_n1672_48),
    .I2(u_usb_device_controller_usb_control_inst_n1672_49) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s41 .INIT=8'h10;
  LUT4 \u_usb_device_controller/usb_control_inst/n1672_s42  (
    .F(u_usb_device_controller_usb_control_inst_n1672_46),
    .I0(u_usb_device_controller_usb_control_inst_n1649_23),
    .I1(u_usb_device_controller_usb_control_inst_n1661_17),
    .I2(u_usb_device_controller_usb_control_inst_n1678_42),
    .I3(u_usb_device_controller_usb_control_inst_n1678_40) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s42 .INIT=16'hB0BB;
  LUT2 \u_usb_device_controller/usb_control_inst/n1678_s38  (
    .F(u_usb_device_controller_usb_control_inst_n1678_42),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1678_s38 .INIT=4'h1;
  LUT3 \u_usb_device_controller/usb_control_inst/n1678_s39  (
    .F(u_usb_device_controller_usb_control_inst_n1678_43),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1678_s39 .INIT=8'h0B;
  LUT4 \u_usb_device_controller/usb_control_inst/n1678_s40  (
    .F(u_usb_device_controller_usb_control_inst_n1678_44),
    .I0(u_usb_device_controller_usb_control_inst_s_test_sel),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I3(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1678_s40 .INIT=16'hC0BF;
  LUT4 \u_usb_device_controller/usb_control_inst/n1680_s42  (
    .F(u_usb_device_controller_usb_control_inst_n1680_46),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I3(u_usb_device_controller_usb_control_inst_n1680_48) 
);
defparam \u_usb_device_controller/usb_control_inst/n1680_s42 .INIT=16'h4532;
  LUT4 \u_usb_device_controller/usb_control_inst/n1680_s43  (
    .F(u_usb_device_controller_usb_control_inst_n1680_47),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I3(u_usb_device_controller_usb_control_inst_n1678_44) 
);
defparam \u_usb_device_controller/usb_control_inst/n1680_s43 .INIT=16'h4532;
  LUT3 \u_usb_device_controller/usb_control_inst/n1684_s37  (
    .F(u_usb_device_controller_usb_control_inst_n1684_41),
    .I0(u_usb_device_controller_usb_control_inst_s_state[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[1]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1684_s37 .INIT=8'h10;
  LUT2 \u_usb_device_controller/usb_control_inst/n1684_s38  (
    .F(u_usb_device_controller_usb_control_inst_n1684_42),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1684_s38 .INIT=4'h1;
  LUT4 \u_usb_device_controller/usb_control_inst/n1686_s37  (
    .F(u_usb_device_controller_usb_control_inst_n1686_41),
    .I0(u_usb_device_controller_usb_control_inst_n1686_43),
    .I1(u_usb_device_controller_usb_control_inst_n1686_44),
    .I2(u_usb_device_controller_usb_control_inst_n1686_50),
    .I3(u_usb_device_controller_usb_control_inst_s_setupptr[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1686_s37 .INIT=16'hF0EE;
  LUT3 \u_usb_device_controller/usb_control_inst/n1686_s38  (
    .F(u_usb_device_controller_usb_control_inst_n1686_42),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .I2(u_usb_device_controller_usb_control_inst_n1684_40) 
);
defparam \u_usb_device_controller/usb_control_inst/n1686_s38 .INIT=8'h07;
  LUT4 \u_usb_device_controller/usb_control_inst/n1690_s33  (
    .F(u_usb_device_controller_usb_control_inst_n1690_37),
    .I0(u_usb_device_controller_usb_control_inst_n1876_9),
    .I1(u_usb_device_controller_usb_control_inst_n435_20),
    .I2(u_usb_device_controller_usb_control_inst_n1690_39),
    .I3(u_usb_device_controller_usb_control_inst_n1629) 
);
defparam \u_usb_device_controller/usb_control_inst/n1690_s33 .INIT=16'h0700;
  LUT2 \u_usb_device_controller/usb_control_inst/n1690_s34  (
    .F(u_usb_device_controller_usb_control_inst_n1690_38),
    .I0(u_usb_device_controller_usb_control_inst_s_test_sel),
    .I1(u_usb_device_controller_usb_control_inst_n2902_5) 
);
defparam \u_usb_device_controller/usb_control_inst/n1690_s34 .INIT=4'h4;
  LUT2 \u_usb_device_controller/usb_control_inst/n1709_s13  (
    .F(u_usb_device_controller_usb_control_inst_n1709_17),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1709_s13 .INIT=4'h4;
  LUT2 \u_usb_device_controller/usb_control_inst/n1649_s15  (
    .F(u_usb_device_controller_usb_control_inst_n1649_19),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[4]),
    .I1(u_usb_device_controller_usb_control_inst_n1652_24) 
);
defparam \u_usb_device_controller/usb_control_inst/n1649_s15 .INIT=4'h8;
  LUT4 \u_usb_device_controller/usb_control_inst/n1649_s17  (
    .F(u_usb_device_controller_usb_control_inst_n1649_21),
    .I0(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[7]),
    .I3(u_usb_device_controller_usb_control_inst_s_state[8]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1649_s17 .INIT=16'h0110;
  LUT4 \u_usb_device_controller/usb_control_inst/n1652_s15  (
    .F(u_usb_device_controller_usb_control_inst_n1652_19),
    .I0(u_usb_device_controller_usb_control_inst_s_state[7]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I3(u_usb_device_controller_usb_control_inst_s_state[8]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1652_s15 .INIT=16'h0110;
  LUT2 \u_usb_device_controller/u_usb_packet/n626_s40  (
    .F(u_usb_device_controller_u_usb_packet_n626_44),
    .I0(txval_i_d),
    .I1(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/u_usb_packet/n626_s40 .INIT=4'h4;
  LUT2 \u_usb_device_controller/u_usb_packet/n626_s41  (
    .F(u_usb_device_controller_u_usb_packet_n626_45),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(u_usb_device_controller_n1615_15) 
);
defparam \u_usb_device_controller/u_usb_packet/n626_s41 .INIT=4'h1;
  LUT2 \u_usb_device_controller/u_usb_packet/n626_s42  (
    .F(u_usb_device_controller_u_usb_packet_n626_46),
    .I0(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I1(u_usb_device_controller_u_usb_init_usbp_chirpk) 
);
defparam \u_usb_device_controller/u_usb_packet/n626_s42 .INIT=4'h1;
  LUT2 \u_usb_device_controller/u_usb_packet/n628_s44  (
    .F(u_usb_device_controller_u_usb_packet_n628_48),
    .I0(u_usb_device_controller_u_usb_packet_n628_49),
    .I1(u_usb_device_controller_u_usb_packet_n628_50) 
);
defparam \u_usb_device_controller/u_usb_packet/n628_s44 .INIT=4'h8;
  LUT4 \u_usb_device_controller/u_usb_packet/n633_s36  (
    .F(u_usb_device_controller_u_usb_packet_n633_40),
    .I0(u_usb_device_controller_u_usb_packet_n615_44),
    .I1(u_usb_device_controller_u_usb_packet_s_state_11_22),
    .I2(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I3(u_usb_device_controller_u_usb_packet_s_rxerror) 
);
defparam \u_usb_device_controller/u_usb_packet/n633_s36 .INIT=16'hE000;
  LUT4 \u_usb_device_controller/u_usb_packet/n633_s37  (
    .F(u_usb_device_controller_u_usb_packet_n633_41),
    .I0(u_usb_device_controller_u_usb_packet_n628_48),
    .I1(u_usb_device_controller_u_usb_packet_s_state_11_22),
    .I2(u_usb_device_controller_u_usb_packet_n633_43),
    .I3(u_usb_device_controller_usb_transact_inst_n1565_4) 
);
defparam \u_usb_device_controller/u_usb_packet/n633_s37 .INIT=16'hF400;
  LUT3 \u_usb_device_controller/u_usb_packet/n633_s38  (
    .F(u_usb_device_controller_u_usb_packet_n633_42),
    .I0(u_usb_device_controller_u_usb_packet_n633_44),
    .I1(u_usb_device_controller_u_usb_packet_s_txready),
    .I2(u_usb_device_controller_u_usb_packet_n920_6) 
);
defparam \u_usb_device_controller/u_usb_packet/n633_s38 .INIT=8'hCA;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1091_s47  (
    .F(u_usb_device_controller_usb_transact_inst_n1091_52),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[9]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[8]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1091_s47 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1095_s43  (
    .F(u_usb_device_controller_usb_transact_inst_n1095_47),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[5]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[7]),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[6]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1095_s43 .INIT=16'h0100;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1101_s41  (
    .F(u_usb_device_controller_usb_transact_inst_n1101_45),
    .I0(u_usb_device_controller_usb_transact_inst_s_ping),
    .I1(u_usb_device_controller_usb_transact_inst_s_in) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1101_s41 .INIT=4'h1;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1109_s45  (
    .F(u_usb_device_controller_usb_transact_inst_n1109_49),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_usb_transact_inst_n1111_18),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I3(u_usb_device_controller_u_usb_packet_s_rxvalid) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1109_s45 .INIT=16'hF100;
  LUT2 \u_usb_device_controller/usb_transact_inst/n1138_s26  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_31),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[7]),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[8]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s26 .INIT=4'h1;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1072_s16  (
    .F(u_usb_device_controller_usb_transact_inst_n1072_22),
    .I0(u_usb_device_controller_u_usb_packet_n784_20),
    .I1(u_usb_device_controller_u_usb_packet_n622_46),
    .I2(u_usb_device_controller_u_usb_packet_n800_6) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1072_s16 .INIT=8'h0B;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1159_s22  (
    .F(u_usb_device_controller_usb_transact_inst_n1159_27),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid_3_16),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_s_nyet) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1159_s22 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/usb_control_inst/n1860_s26  (
    .F(u_usb_device_controller_usb_control_inst_n1860_31),
    .I0(u_usb_device_controller_usb_control_inst_n1860_33),
    .I1(u_usb_device_controller_usb_control_inst_n645_45),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1860_s26 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usb_control_inst/n1860_s27  (
    .F(u_usb_device_controller_usb_control_inst_n1860_32),
    .I0(u_usb_device_controller_usb_control_inst_online_o_d),
    .I1(inf_alter_i_d[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1860_s27 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/usb_control_inst/s_ctlparam_7_s5  (
    .F(u_usb_device_controller_usb_control_inst_s_ctlparam_7_8),
    .I0(u_usb_device_controller_usb_control_inst_s_test_sel),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I2(u_usb_device_controller_usb_control_inst_n2902_5),
    .I3(u_usb_device_controller_usb_control_inst_s_setupptr[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/s_ctlparam_7_s5 .INIT=16'h7F00;
  LUT2 \u_usb_device_controller/test_packet_inst/cnt_11_s6  (
    .F(u_usb_device_controller_test_packet_inst_cnt_11_11),
    .I0(u_usb_device_controller_test_packet_inst_cnt[4]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[5]) 
);
defparam \u_usb_device_controller/test_packet_inst/cnt_11_s6 .INIT=4'h8;
  LUT3 \u_usb_device_controller/test_packet_inst/cnt_11_s7  (
    .F(u_usb_device_controller_test_packet_inst_cnt_11_12),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[1]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_testmode[6]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_testmode[7]) 
);
defparam \u_usb_device_controller/test_packet_inst/cnt_11_s7 .INIT=8'h01;
  LUT4 \u_usb_device_controller/test_packet_inst/cnt_11_s8  (
    .F(u_usb_device_controller_test_packet_inst_cnt_11_13),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_testmode[4]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_testmode[5]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_testmode[2]) 
);
defparam \u_usb_device_controller/test_packet_inst/cnt_11_s8 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/test_packet_inst/test_data_6_s6  (
    .F(u_usb_device_controller_test_packet_inst_test_data_6_9),
    .I0(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[2]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[3]) 
);
defparam \u_usb_device_controller/test_packet_inst/test_data_6_s6 .INIT=16'h001F;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_2_s11  (
    .F(u_usb_device_controller_u_usb_init_s_state_2_16),
    .I0(u_usb_device_controller_u_usb_init_s_linestate[1]),
    .I1(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I2(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .I3(u_usb_device_controller_u_usb_init_n414) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_2_s11 .INIT=16'hD000;
  LUT2 \u_usb_device_controller/test_packet_inst/n318_s7  (
    .F(u_usb_device_controller_test_packet_inst_n318_11),
    .I0(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[2]) 
);
defparam \u_usb_device_controller/test_packet_inst/n318_s7 .INIT=4'h1;
  LUT4 \u_usb_device_controller/test_packet_inst/n318_s8  (
    .F(u_usb_device_controller_test_packet_inst_n318_12),
    .I0(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[4]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[2]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[3]) 
);
defparam \u_usb_device_controller/test_packet_inst/n318_s8 .INIT=16'h233F;
  LUT4 \u_usb_device_controller/test_packet_inst/n318_s9  (
    .F(u_usb_device_controller_test_packet_inst_n318_13),
    .I0(u_usb_device_controller_test_packet_inst_cnt[8]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[9]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[10]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[11]) 
);
defparam \u_usb_device_controller/test_packet_inst/n318_s9 .INIT=16'h0001;
  LUT2 \u_usb_device_controller/test_packet_inst/n318_s10  (
    .F(u_usb_device_controller_test_packet_inst_n318_14),
    .I0(u_usb_device_controller_test_packet_inst_cnt[4]),
    .I1(u_usb_device_controller_test_packet_inst_n312_13) 
);
defparam \u_usb_device_controller/test_packet_inst/n318_s10 .INIT=4'h4;
  LUT4 \u_usb_device_controller/test_packet_inst/n317_s7  (
    .F(u_usb_device_controller_test_packet_inst_n317_11),
    .I0(u_usb_device_controller_test_packet_inst_cnt_11_11),
    .I1(u_usb_device_controller_test_packet_inst_cnt[2]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[0]) 
);
defparam \u_usb_device_controller/test_packet_inst/n317_s7 .INIT=16'h4FFB;
  LUT4 \u_usb_device_controller/test_packet_inst/n311_s6  (
    .F(u_usb_device_controller_test_packet_inst_n311_10),
    .I0(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[4]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[2]) 
);
defparam \u_usb_device_controller/test_packet_inst/n311_s6 .INIT=16'h1400;
  LUT4 \u_usb_device_controller/u_usb_init/n219_s21  (
    .F(u_usb_device_controller_u_usb_init_n219_29),
    .I0(u_usb_device_controller_u_usb_init_s_chirpcnt_2_9),
    .I1(u_usb_device_controller_u_usb_init_n212_43),
    .I2(u_usb_device_controller_u_usb_init_n219_30),
    .I3(u_usb_device_controller_u_usb_init_s_state_0_4) 
);
defparam \u_usb_device_controller/u_usb_init/n219_s21 .INIT=16'h00FE;
  LUT2 \u_usb_device_controller/n1534_s23  (
    .F(u_usb_device_controller_n1534_30),
    .I0(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I1(u_usb_device_controller_usb_transact_inst_s_in_valid) 
);
defparam \u_usb_device_controller/n1534_s23 .INIT=4'h4;
  LUT4 \u_usb_device_controller/n1534_s24  (
    .F(u_usb_device_controller_n1534_31),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I1(u_usb_device_controller_cur_state[0]),
    .I2(u_usb_device_controller_cur_state[1]),
    .I3(u_usb_device_controller_rxact_o_d_3) 
);
defparam \u_usb_device_controller/n1534_s24 .INIT=16'h0700;
  LUT4 \u_usb_device_controller/n1534_s25  (
    .F(u_usb_device_controller_n1534_32),
    .I0(u_usb_device_controller_n1534_35),
    .I1(u_usb_device_controller_n1534_30),
    .I2(u_usb_device_controller_cur_state[0]),
    .I3(u_usb_device_controller_rxdat_d0_7_9) 
);
defparam \u_usb_device_controller/n1534_s25 .INIT=16'h0007;
  LUT4 \u_usb_device_controller/n1534_s26  (
    .F(u_usb_device_controller_n1534_33),
    .I0(u_usb_device_controller_n1465_3),
    .I1(u_usb_device_controller_cur_state[0]),
    .I2(u_usb_device_controller_n1534_30),
    .I3(u_usb_device_controller_cur_state[1]) 
);
defparam \u_usb_device_controller/n1534_s26 .INIT=16'hBF00;
  LUT4 \u_usb_device_controller/n1534_s27  (
    .F(u_usb_device_controller_n1534_34),
    .I0(u_usb_device_controller_s_halt_out),
    .I1(u_usb_device_controller_s_endpt_rxrdy),
    .I2(u_usb_device_controller_setup_o_d_3),
    .I3(u_usb_device_controller_rxdat_d0_7_9) 
);
defparam \u_usb_device_controller/n1534_s27 .INIT=16'h4000;
  LUT2 \u_usb_device_controller/n1529_s22  (
    .F(u_usb_device_controller_n1529_28),
    .I0(u_usb_device_controller_s_endpt_rxrdy),
    .I1(u_usb_device_controller_usb_transact_inst_T_PING_2) 
);
defparam \u_usb_device_controller/n1529_s22 .INIT=4'h4;
  LUT4 \u_usb_device_controller/n1529_s23  (
    .F(u_usb_device_controller_n1529_29),
    .I0(u_usb_device_controller_usb_transact_inst_s_setup_2),
    .I1(u_usb_device_controller_usb_transact_inst_s_out_valid),
    .I2(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/n1529_s23 .INIT=16'hF100;
  LUT2 \u_usb_device_controller/usbc_dsclen_0_s11  (
    .F(u_usb_device_controller_usbc_dsclen_0_16),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s11 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usbc_dsclen_0_s12  (
    .F(u_usb_device_controller_usbc_dsclen_0_17),
    .I0(desc_have_strings_i_d),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s12 .INIT=16'hF08C;
  LUT4 \u_usb_device_controller/usbc_dsclen_0_s13  (
    .F(u_usb_device_controller_usbc_dsclen_0_18),
    .I0(u_usb_device_controller_usbc_dsclen_0_20),
    .I1(u_usb_device_controller_usbc_dsclen_1_24),
    .I2(u_usb_device_controller_usbc_dsclen_0_21),
    .I3(u_usb_device_controller_usbc_dsclen_0_22) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s13 .INIT=16'h00BF;
  LUT4 \u_usb_device_controller/usbc_dsclen_0_s14  (
    .F(u_usb_device_controller_usbc_dsclen_0_19),
    .I0(u_usb_device_controller_usbc_dsclen_0_23),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_len_i_d[0]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s14 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/usbc_dsclen_1_s11  (
    .F(u_usb_device_controller_usbc_dsclen_1_16),
    .I0(desc_hscfg_len_i_d[1]),
    .I1(desc_fscfg_len_i_d[1]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usb_control_inst_n1836_10) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s11 .INIT=16'hCA00;
  LUT4 \u_usb_device_controller/usbc_dsclen_1_s13  (
    .F(u_usb_device_controller_usbc_dsclen_1_18),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(desc_strproduct_len_i_d[1]),
    .I2(desc_strserial_len_i_d[1]),
    .I3(u_usb_device_controller_usb_control_inst_n1705_16) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s13 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/usbc_dsclen_1_s15  (
    .F(u_usb_device_controller_usbc_dsclen_1_20),
    .I0(desc_dev_len_i_d[1]),
    .I1(u_usb_device_controller_usbc_dsclen_1_22),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s15 .INIT=16'h0305;
  LUT4 \u_usb_device_controller/usbc_dsclen_2_s11  (
    .F(u_usb_device_controller_usbc_dsclen_2_16),
    .I0(u_usb_device_controller_usbc_dsclen_2_18),
    .I1(u_usb_device_controller_usbc_dsclen_2_19),
    .I2(u_usb_device_controller_usbc_dsclen_2_20),
    .I3(u_usb_device_controller_usb_control_inst_n1836_9) 
);
defparam \u_usb_device_controller/usbc_dsclen_2_s11 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/usbc_dsclen_2_s12  (
    .F(u_usb_device_controller_usbc_dsclen_2_17),
    .I0(desc_hscfg_len_i_d[2]),
    .I1(desc_fscfg_len_i_d[2]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_2_s12 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/usbc_dsclen_3_s10  (
    .F(u_usb_device_controller_usbc_dsclen_3_15),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(desc_strvendor_len_i_d[3]),
    .I2(u_usb_device_controller_usbc_dsclen_3_18),
    .I3(u_usb_device_controller_usbc_dsclen_1_24) 
);
defparam \u_usb_device_controller/usbc_dsclen_3_s10 .INIT=16'h8F00;
  LUT3 \u_usb_device_controller/usbc_dsclen_3_s11  (
    .F(u_usb_device_controller_usbc_dsclen_3_16),
    .I0(desc_dev_len_i_d[3]),
    .I1(u_usb_device_controller_usbc_dsclen_3_19),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_3_s11 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/usbc_dsclen_3_s12  (
    .F(u_usb_device_controller_usbc_dsclen_3_17),
    .I0(u_usb_device_controller_usbc_dsclen_3_20),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_len_i_d[3]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/usbc_dsclen_3_s12 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/usbc_dsclen_4_s11  (
    .F(u_usb_device_controller_usbc_dsclen_4_16),
    .I0(desc_fscfg_len_i_d[4]),
    .I1(desc_hscfg_len_i_d[4]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I3(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_4_s11 .INIT=16'h0C0A;
  LUT4 \u_usb_device_controller/usbc_dsclen_4_s12  (
    .F(u_usb_device_controller_usbc_dsclen_4_17),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(desc_strvendor_len_i_d[4]),
    .I2(u_usb_device_controller_usbc_dsclen_4_19),
    .I3(u_usb_device_controller_usbc_dsclen_1_24) 
);
defparam \u_usb_device_controller/usbc_dsclen_4_s12 .INIT=16'h8F00;
  LUT3 \u_usb_device_controller/usbc_dsclen_4_s13  (
    .F(u_usb_device_controller_usbc_dsclen_4_18),
    .I0(desc_hscfg_len_i_d[4]),
    .I1(desc_fscfg_len_i_d[4]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_4_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/usbc_dsclen_5_s10  (
    .F(u_usb_device_controller_usbc_dsclen_5_15),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(desc_strvendor_len_i_d[5]),
    .I2(u_usb_device_controller_usbc_dsclen_5_18),
    .I3(u_usb_device_controller_usbc_dsclen_1_24) 
);
defparam \u_usb_device_controller/usbc_dsclen_5_s10 .INIT=16'h8F00;
  LUT4 \u_usb_device_controller/usbc_dsclen_5_s11  (
    .F(u_usb_device_controller_usbc_dsclen_5_16),
    .I0(u_usb_device_controller_usbc_dsclen_5_19),
    .I1(u_usb_device_controller_usbc_dsclen_0_16),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I3(desc_dev_len_i_d[5]) 
);
defparam \u_usb_device_controller/usbc_dsclen_5_s11 .INIT=16'h7077;
  LUT4 \u_usb_device_controller/usbc_dsclen_5_s12  (
    .F(u_usb_device_controller_usbc_dsclen_5_17),
    .I0(u_usb_device_controller_usbc_dsclen_5_20),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_len_i_d[5]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/usbc_dsclen_5_s12 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/usbc_dsclen_6_s11  (
    .F(u_usb_device_controller_usbc_dsclen_6_16),
    .I0(u_usb_device_controller_usbc_dsclen_6_18),
    .I1(u_usb_device_controller_usbc_dsclen_1_24),
    .I2(u_usb_device_controller_usbc_dsclen_6_19),
    .I3(u_usb_device_controller_usbc_dsclen_6_20) 
);
defparam \u_usb_device_controller/usbc_dsclen_6_s11 .INIT=16'h00BF;
  LUT4 \u_usb_device_controller/usbc_dsclen_6_s12  (
    .F(u_usb_device_controller_usbc_dsclen_6_17),
    .I0(desc_hscfg_len_i_d[6]),
    .I1(desc_fscfg_len_i_d[6]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usb_control_inst_n1836_10) 
);
defparam \u_usb_device_controller/usbc_dsclen_6_s12 .INIT=16'hCA00;
  LUT4 \u_usb_device_controller/usbc_dsclen_7_s10  (
    .F(u_usb_device_controller_usbc_dsclen_7_15),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(desc_strvendor_len_i_d[7]),
    .I2(u_usb_device_controller_usbc_dsclen_7_18),
    .I3(u_usb_device_controller_usbc_dsclen_1_24) 
);
defparam \u_usb_device_controller/usbc_dsclen_7_s10 .INIT=16'h8F00;
  LUT4 \u_usb_device_controller/usbc_dsclen_7_s11  (
    .F(u_usb_device_controller_usbc_dsclen_7_16),
    .I0(u_usb_device_controller_usbc_dsclen_7_19),
    .I1(u_usb_device_controller_usbc_dsclen_0_16),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I3(desc_dev_len_i_d[7]) 
);
defparam \u_usb_device_controller/usbc_dsclen_7_s11 .INIT=16'h7077;
  LUT4 \u_usb_device_controller/usbc_dsclen_7_s12  (
    .F(u_usb_device_controller_usbc_dsclen_7_17),
    .I0(u_usb_device_controller_usbc_dsclen_7_20),
    .I1(u_usb_device_controller_usb_control_inst_n1836_10),
    .I2(desc_qual_len_i_d[7]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]) 
);
defparam \u_usb_device_controller/usbc_dsclen_7_s12 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/descrom_start_0_s11  (
    .F(u_usb_device_controller_descrom_start_0_16),
    .I0(desc_fscfg_addr_i_d[0]),
    .I1(desc_hscfg_addr_i_d[0]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_0_s11 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/descrom_start_0_s12  (
    .F(u_usb_device_controller_descrom_start_0_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[0]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_0_19) 
);
defparam \u_usb_device_controller/descrom_start_0_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_0_s13  (
    .F(u_usb_device_controller_descrom_start_0_18),
    .I0(desc_hscfg_addr_i_d[0]),
    .I1(desc_fscfg_addr_i_d[0]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_0_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_1_s11  (
    .F(u_usb_device_controller_descrom_start_1_16),
    .I0(desc_fscfg_addr_i_d[1]),
    .I1(desc_hscfg_addr_i_d[1]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_1_s11 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/descrom_start_1_s12  (
    .F(u_usb_device_controller_descrom_start_1_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[1]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_1_19) 
);
defparam \u_usb_device_controller/descrom_start_1_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_1_s13  (
    .F(u_usb_device_controller_descrom_start_1_18),
    .I0(desc_hscfg_addr_i_d[1]),
    .I1(desc_fscfg_addr_i_d[1]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_1_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_2_s11  (
    .F(u_usb_device_controller_descrom_start_2_16),
    .I0(desc_fscfg_addr_i_d[2]),
    .I1(desc_hscfg_addr_i_d[2]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_2_s11 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/descrom_start_2_s12  (
    .F(u_usb_device_controller_descrom_start_2_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[2]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_2_19) 
);
defparam \u_usb_device_controller/descrom_start_2_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_2_s13  (
    .F(u_usb_device_controller_descrom_start_2_18),
    .I0(desc_hscfg_addr_i_d[2]),
    .I1(desc_fscfg_addr_i_d[2]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_2_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_3_s11  (
    .F(u_usb_device_controller_descrom_start_3_16),
    .I0(desc_fscfg_addr_i_d[3]),
    .I1(desc_hscfg_addr_i_d[3]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_3_s11 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/descrom_start_3_s12  (
    .F(u_usb_device_controller_descrom_start_3_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[3]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_3_19) 
);
defparam \u_usb_device_controller/descrom_start_3_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_3_s13  (
    .F(u_usb_device_controller_descrom_start_3_18),
    .I0(desc_hscfg_addr_i_d[3]),
    .I1(desc_fscfg_addr_i_d[3]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_3_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_4_s11  (
    .F(u_usb_device_controller_descrom_start_4_16),
    .I0(desc_fscfg_addr_i_d[4]),
    .I1(desc_hscfg_addr_i_d[4]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_4_s11 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/descrom_start_4_s12  (
    .F(u_usb_device_controller_descrom_start_4_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[4]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_4_19) 
);
defparam \u_usb_device_controller/descrom_start_4_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_4_s13  (
    .F(u_usb_device_controller_descrom_start_4_18),
    .I0(desc_hscfg_addr_i_d[4]),
    .I1(desc_fscfg_addr_i_d[4]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_4_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_5_s11  (
    .F(u_usb_device_controller_descrom_start_5_16),
    .I0(desc_fscfg_addr_i_d[5]),
    .I1(desc_hscfg_addr_i_d[5]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_5_s11 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/descrom_start_5_s12  (
    .F(u_usb_device_controller_descrom_start_5_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[5]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_5_19) 
);
defparam \u_usb_device_controller/descrom_start_5_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_5_s13  (
    .F(u_usb_device_controller_descrom_start_5_18),
    .I0(desc_hscfg_addr_i_d[5]),
    .I1(desc_fscfg_addr_i_d[5]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_5_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_6_s11  (
    .F(u_usb_device_controller_descrom_start_6_16),
    .I0(desc_fscfg_addr_i_d[6]),
    .I1(desc_hscfg_addr_i_d[6]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_6_s11 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/descrom_start_6_s12  (
    .F(u_usb_device_controller_descrom_start_6_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[6]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_6_19) 
);
defparam \u_usb_device_controller/descrom_start_6_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_6_s13  (
    .F(u_usb_device_controller_descrom_start_6_18),
    .I0(desc_hscfg_addr_i_d[6]),
    .I1(desc_fscfg_addr_i_d[6]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_6_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_7_s11  (
    .F(u_usb_device_controller_descrom_start_7_16),
    .I0(desc_fscfg_addr_i_d[7]),
    .I1(desc_hscfg_addr_i_d[7]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_7_s11 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/descrom_start_7_s12  (
    .F(u_usb_device_controller_descrom_start_7_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[7]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_7_19) 
);
defparam \u_usb_device_controller/descrom_start_7_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_7_s13  (
    .F(u_usb_device_controller_descrom_start_7_18),
    .I0(desc_hscfg_addr_i_d[7]),
    .I1(desc_fscfg_addr_i_d[7]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_7_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_8_s11  (
    .F(u_usb_device_controller_descrom_start_8_16),
    .I0(desc_fscfg_addr_i_d[8]),
    .I1(desc_hscfg_addr_i_d[8]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_8_s11 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/descrom_start_8_s12  (
    .F(u_usb_device_controller_descrom_start_8_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[8]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_8_19) 
);
defparam \u_usb_device_controller/descrom_start_8_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_8_s13  (
    .F(u_usb_device_controller_descrom_start_8_18),
    .I0(desc_hscfg_addr_i_d[8]),
    .I1(desc_fscfg_addr_i_d[8]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_8_s13 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_9_s11  (
    .F(u_usb_device_controller_descrom_start_9_16),
    .I0(desc_hscfg_addr_i_d[9]),
    .I1(desc_fscfg_addr_i_d[9]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usbc_dsclen_0_16) 
);
defparam \u_usb_device_controller/descrom_start_9_s11 .INIT=16'h5300;
  LUT4 \u_usb_device_controller/descrom_start_9_s12  (
    .F(u_usb_device_controller_descrom_start_9_17),
    .I0(u_usb_device_controller_usb_control_inst_n1836_13),
    .I1(desc_strproduct_addr_i_d[9]),
    .I2(u_usb_device_controller_usbc_dsclen_1_21),
    .I3(u_usb_device_controller_descrom_start_9_19) 
);
defparam \u_usb_device_controller/descrom_start_9_s12 .INIT=16'h7000;
  LUT3 \u_usb_device_controller/descrom_start_9_s13  (
    .F(u_usb_device_controller_descrom_start_9_18),
    .I0(desc_hscfg_addr_i_d[9]),
    .I1(desc_fscfg_addr_i_d[9]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/descrom_start_9_s13 .INIT=8'hCA;
  LUT2 \u_usb_device_controller/usb_transact_inst/txpop_o_d_s3  (
    .F(u_usb_device_controller_usb_transact_inst_txpop_o_d_7),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[9]) 
);
defparam \u_usb_device_controller/usb_transact_inst/txpop_o_d_s3 .INIT=4'h4;
  LUT4 \u_usb_device_controller/test_packet_inst/n313_s5  (
    .F(u_usb_device_controller_test_packet_inst_n313_9),
    .I0(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[2]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[4]) 
);
defparam \u_usb_device_controller/test_packet_inst/n313_s5 .INIT=16'hBFC8;
  LUT3 \u_usb_device_controller/u_usb_packet/n774_s4  (
    .F(u_usb_device_controller_u_usb_packet_n774_8),
    .I0(u_usb_device_controller_u_usb_packet_n919_5),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[2]),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54) 
);
defparam \u_usb_device_controller/u_usb_packet/n774_s4 .INIT=8'hB0;
  LUT2 \u_usb_device_controller/u_usb_packet/n774_s5  (
    .F(u_usb_device_controller_u_usb_packet_n774_9),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]),
    .I1(u_usb_device_controller_u_usb_packet_n912_14) 
);
defparam \u_usb_device_controller/u_usb_packet/n774_s5 .INIT=4'h8;
  LUT3 \u_usb_device_controller/u_usb_packet/n774_s6  (
    .F(u_usb_device_controller_u_usb_packet_n774_10),
    .I0(u_usb_device_controller_u_usb_packet_n919_5),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[3]),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54) 
);
defparam \u_usb_device_controller/u_usb_packet/n774_s6 .INIT=8'hB0;
  LUT2 \u_usb_device_controller/u_usb_packet/n774_s7  (
    .F(u_usb_device_controller_u_usb_packet_n774_11),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .I1(u_usb_device_controller_u_usb_packet_n912_14) 
);
defparam \u_usb_device_controller/u_usb_packet/n774_s7 .INIT=4'h8;
  LUT3 \u_usb_device_controller/u_usb_packet/n771_s4  (
    .F(u_usb_device_controller_u_usb_packet_n771_8),
    .I0(u_usb_device_controller_u_usb_packet_n919_5),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[0]),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s4 .INIT=8'hB0;
  LUT2 \u_usb_device_controller/u_usb_packet/n771_s5  (
    .F(u_usb_device_controller_u_usb_packet_n771_9),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .I1(u_usb_device_controller_u_usb_packet_n912_14) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s5 .INIT=4'h8;
  LUT3 \u_usb_device_controller/u_usb_packet/n771_s6  (
    .F(u_usb_device_controller_u_usb_packet_n771_10),
    .I0(u_usb_device_controller_u_usb_packet_n771_13),
    .I1(u_usb_device_controller_u_usb_packet_n328_12),
    .I2(u_usb_device_controller_u_usb_packet_n771_14) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s6 .INIT=8'hD0;
  LUT3 \u_usb_device_controller/u_usb_packet/n771_s7  (
    .F(u_usb_device_controller_u_usb_packet_n771_11),
    .I0(u_usb_device_controller_u_usb_packet_n626_42),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[3]),
    .I2(u_usb_device_controller_u_usb_packet_n622_46) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s7 .INIT=8'hE0;
  LUT2 \u_usb_device_controller/u_usb_packet/n771_s8  (
    .F(u_usb_device_controller_u_usb_packet_n771_12),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I1(u_usb_device_controller_u_usb_packet_crc16_buf_15_14) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s8 .INIT=4'h8;
  LUT4 \u_usb_device_controller/u_usb_packet/n767_s4  (
    .F(u_usb_device_controller_u_usb_packet_n767_8),
    .I0(u_usb_device_controller_u_usb_packet_n328_24),
    .I1(u_usb_device_controller_u_usb_packet_n919_5),
    .I2(u_usb_device_controller_u_usb_packet_n767_9),
    .I3(u_usb_device_controller_u_usb_packet_n767_10) 
);
defparam \u_usb_device_controller/u_usb_packet/n767_s4 .INIT=16'h004F;
  LUT2 \u_usb_device_controller/u_usb_packet/crc5_buf_4_s7  (
    .F(u_usb_device_controller_u_usb_packet_crc5_buf_4_11),
    .I0(u_usb_device_controller_u_usb_packet_s_rxerror),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact) 
);
defparam \u_usb_device_controller/u_usb_packet/crc5_buf_4_s7 .INIT=4'h4;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1133_s21  (
    .F(u_usb_device_controller_usb_transact_inst_n1133_27),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[4]),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[5]),
    .I2(u_usb_device_controller_usb_transact_inst_wait_count[6]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1133_s21 .INIT=8'h01;
  LUT2 \u_usb_device_controller/u_usb_packet/n579_s15  (
    .F(u_usb_device_controller_u_usb_packet_n579_21),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf[2]) 
);
defparam \u_usb_device_controller/u_usb_packet/n579_s15 .INIT=4'h6;
  LUT3 \u_usb_device_controller/u_usb_packet/n579_s16  (
    .F(u_usb_device_controller_u_usb_packet_n579_22),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .I1(u_usb_device_controller_u_usb_packet_crc5_buf[0]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]) 
);
defparam \u_usb_device_controller/u_usb_packet/n579_s16 .INIT=8'h96;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_7_s4  (
    .F(u_usb_device_controller_utmi_dataout_o_d_7_8),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_testmode[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_testmode[4]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_testmode[5]) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_7_s4 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/n2024_s4  (
    .F(u_usb_device_controller_n2024_7),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscoff[4]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscoff[5]) 
);
defparam \u_usb_device_controller/n2024_s4 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/u_usb_packet/n784_s10  (
    .F(u_usb_device_controller_u_usb_packet_n784_13),
    .I0(u_usb_device_controller_u_usb_packet_n626_42),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[1]),
    .I2(u_usb_device_controller_u_usb_packet_n919_5),
    .I3(u_usb_device_controller_usb_transact_inst_n1091_54) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s10 .INIT=16'hAC00;
  LUT4 \u_usb_device_controller/u_usb_packet/n785_s5  (
    .F(u_usb_device_controller_u_usb_packet_n785_8),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[7]),
    .I1(u_usb_device_controller_u_usb_packet_n620),
    .I2(u_usb_device_controller_u_usb_packet_s_dataout[0]),
    .I3(u_usb_device_controller_u_usb_packet_n782_8) 
);
defparam \u_usb_device_controller/u_usb_packet/n785_s5 .INIT=16'h0BBB;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s11  (
    .F(u_usb_device_controller_u_usb_packet_n912_14),
    .I0(u_usb_device_controller_u_usb_packet_s_state[2]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[3]),
    .I2(u_usb_device_controller_u_usb_packet_n784_9),
    .I3(u_usb_device_controller_u_usb_packet_n784_11) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s11 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s12  (
    .F(u_usb_device_controller_u_usb_packet_n912_15),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[5]),
    .I1(u_usb_device_controller_u_usb_packet_crc16_buf[6]),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf[7]),
    .I3(u_usb_device_controller_u_usb_packet_n912_22) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s12 .INIT=16'h0100;
  LUT3 \u_usb_device_controller/u_usb_packet/n912_s13  (
    .F(u_usb_device_controller_u_usb_packet_n912_16),
    .I0(u_usb_device_controller_u_usb_packet_n919_5),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[1]),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s13 .INIT=8'hB0;
  LUT2 \u_usb_device_controller/u_usb_packet/n912_s14  (
    .F(u_usb_device_controller_u_usb_packet_n912_17),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I1(u_usb_device_controller_u_usb_packet_n912_14) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s14 .INIT=4'h8;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s15  (
    .F(u_usb_device_controller_u_usb_packet_n912_18),
    .I0(u_usb_device_controller_u_usb_packet_n575_19),
    .I1(u_usb_device_controller_u_usb_packet_n573_19),
    .I2(u_usb_device_controller_u_usb_packet_n577_19),
    .I3(u_usb_device_controller_u_usb_packet_n577_20) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s15 .INIT=16'hEFF7;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s16  (
    .F(u_usb_device_controller_u_usb_packet_n912_19),
    .I0(u_usb_device_controller_u_usb_packet_s_rxerror),
    .I1(u_usb_device_controller_usb_transact_inst_n1565_4),
    .I2(u_usb_device_controller_u_usb_packet_n579_20),
    .I3(u_usb_device_controller_u_usb_packet_n579_19) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s16 .INIT=16'h0040;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s17  (
    .F(u_usb_device_controller_u_usb_packet_n912_20),
    .I0(u_usb_device_controller_u_usb_packet_n784_11),
    .I1(u_usb_device_controller_u_usb_packet_n920_7),
    .I2(u_usb_device_controller_u_usb_packet_s_state_11_27),
    .I3(u_usb_device_controller_u_usb_packet_n579_20) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s17 .INIT=16'hF077;
  LUT3 \u_usb_device_controller/u_usb_packet/n912_s18  (
    .F(u_usb_device_controller_u_usb_packet_n912_21),
    .I0(u_usb_device_controller_u_usb_packet_n615_42),
    .I1(u_usb_device_controller_u_usb_packet_n615_49),
    .I2(u_usb_device_controller_u_usb_packet_n912_23) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s18 .INIT=8'h0D;
  LUT3 \u_usb_device_controller/usb_control_inst/n2896_s4  (
    .F(u_usb_device_controller_usb_control_inst_n2896_7),
    .I0(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I1(u_usb_device_controller_u_usb_packet_n328_17),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_5_10) 
);
defparam \u_usb_device_controller/usb_control_inst/n2896_s4 .INIT=8'h80;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s33  (
    .F(u_usb_device_controller_u_usb_init_n212_41),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[12]),
    .I1(u_usb_device_controller_u_usb_init_s_timer1[14]),
    .I2(u_usb_device_controller_u_usb_init_s_timer1[15]),
    .I3(u_usb_device_controller_u_usb_init_n212_46) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s33 .INIT=16'h0100;
  LUT3 \u_usb_device_controller/u_usb_init/n212_s34  (
    .F(u_usb_device_controller_u_usb_init_n212_42),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[0]),
    .I1(u_usb_device_controller_u_usb_init_n212_47),
    .I2(u_usb_device_controller_u_usb_init_n212_48) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s34 .INIT=8'h40;
  LUT3 \u_usb_device_controller/u_usb_init/n212_s35  (
    .F(u_usb_device_controller_u_usb_init_n212_43),
    .I0(u_usb_device_controller_u_usb_init_n215_58),
    .I1(u_usb_device_controller_u_usb_init_s_chirpcnt_2_13),
    .I2(u_usb_device_controller_u_usb_init_n212_49) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s35 .INIT=8'h80;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s36  (
    .F(u_usb_device_controller_u_usb_init_n212_44),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[8]),
    .I1(u_usb_device_controller_u_usb_init_s_chirpcnt_2_14),
    .I2(u_usb_device_controller_u_usb_init_n212_50),
    .I3(u_usb_device_controller_u_usb_init_n212_51) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s36 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s37  (
    .F(u_usb_device_controller_u_usb_init_n212_45),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[7]),
    .I1(u_usb_device_controller_u_usb_init_n212_52),
    .I2(u_usb_device_controller_u_usb_init_n212_53),
    .I3(u_usb_device_controller_u_usb_init_n212_54) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s37 .INIT=16'hBF00;
  LUT4 \u_usb_device_controller/u_usb_init/n215_s51  (
    .F(u_usb_device_controller_u_usb_init_n215_58),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[11]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[4]),
    .I2(u_usb_device_controller_u_usb_init_s_state_3_13),
    .I3(u_usb_device_controller_u_usb_init_n215_61) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s51 .INIT=16'h4000;
  LUT3 \u_usb_device_controller/u_usb_init/n215_s52  (
    .F(u_usb_device_controller_u_usb_init_n215_59),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[5]),
    .I1(u_usb_device_controller_u_usb_init_n212_50),
    .I2(u_usb_device_controller_u_usb_init_n215_62) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s52 .INIT=8'h80;
  LUT3 \u_usb_device_controller/u_usb_packet/n328_s16  (
    .F(u_usb_device_controller_u_usb_packet_n328_20),
    .I0(u_usb_device_controller_usb_control_inst_usbc_txdat[1]),
    .I1(txdat_i_d[1]),
    .I2(txval_i_d) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s16 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s17  (
    .F(u_usb_device_controller_u_usb_packet_n328_21),
    .I0(descrom_rdata_i_d[1]),
    .I1(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I2(u_usb_device_controller_u_usb_packet_n328_17),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_5_10) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s17 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s18  (
    .F(u_usb_device_controller_u_usb_packet_n328_22),
    .I0(u_usb_device_controller_usb_transact_inst_n1072_18),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[5]),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_50),
    .I3(u_usb_device_controller_u_usb_packet_n328_25) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s18 .INIT=16'h0007;
  LUT3 \u_usb_device_controller/u_usb_packet/n328_s19  (
    .F(u_usb_device_controller_u_usb_packet_n328_23),
    .I0(u_usb_device_controller_usb_control_inst_usbc_txdat[0]),
    .I1(txdat_i_d[0]),
    .I2(txval_i_d) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s19 .INIT=8'hCA;
  LUT2 \u_usb_device_controller/u_usb_packet/n328_s20  (
    .F(u_usb_device_controller_u_usb_packet_n328_24),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(txdat_i_d[0]) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s20 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usb_control_inst/n1836_s8  (
    .F(u_usb_device_controller_usb_control_inst_n1836_11),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[4]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[5]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[6]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1836_s8 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_3_s8  (
    .F(u_usb_device_controller_u_usb_init_s_state_3_13),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[0]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[1]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[2]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[3]) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s8 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_3_s9  (
    .F(u_usb_device_controller_u_usb_init_s_state_3_14),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[4]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[6]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[14]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[13]) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s9 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s7  (
    .F(u_usb_device_controller_u_usb_init_s_chirpcnt_2_11),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[9]),
    .I1(u_usb_device_controller_u_usb_init_s_timer1[10]),
    .I2(u_usb_device_controller_u_usb_init_s_timer1[13]),
    .I3(u_usb_device_controller_u_usb_init_s_timer1[2]) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s7 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s8  (
    .F(u_usb_device_controller_u_usb_init_s_chirpcnt_2_12),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[4]),
    .I1(u_usb_device_controller_u_usb_init_s_timer1[8]),
    .I2(u_usb_device_controller_u_usb_init_s_timer1[7]),
    .I3(u_usb_device_controller_u_usb_init_s_timer1[5]) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s8 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s9  (
    .F(u_usb_device_controller_u_usb_init_s_chirpcnt_2_13),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[18]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[19]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[8]),
    .I3(u_usb_device_controller_u_usb_init_n212_52) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s9 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s10  (
    .F(u_usb_device_controller_u_usb_init_s_chirpcnt_2_14),
    .I0(u_usb_device_controller_u_usb_init_s_state_3_13),
    .I1(u_usb_device_controller_u_usb_init_n215_61),
    .I2(u_usb_device_controller_u_usb_init_s_state_3_16),
    .I3(u_usb_device_controller_u_usb_init_s_chirpcnt_2_15) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s10 .INIT=16'h8000;
  LUT3 \u_usb_device_controller/u_usb_packet/n615_s43  (
    .F(u_usb_device_controller_u_usb_packet_n615_47),
    .I0(u_usb_device_controller_u_usb_packet_s_state[2]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[3]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[4]) 
);
defparam \u_usb_device_controller/u_usb_packet/n615_s43 .INIT=8'hE9;
  LUT4 \u_usb_device_controller/usb_control_inst/s_answerptr_7_s12  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_7_16),
    .I0(u_usb_device_controller_usb_control_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[5]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I3(u_usb_device_controller_usb_control_inst_n1629_5) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_7_s12 .INIT=16'h0100;
  LUT3 \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s13  (
    .F(u_usb_device_controller_usb_control_inst_s_sendbyte_7_17),
    .I0(u_usb_device_controller_usb_control_inst_n1715_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_n1876_13) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s13 .INIT=8'hD0;
  LUT4 \u_usb_device_controller/u_usb_packet/s_state_11_s20  (
    .F(u_usb_device_controller_u_usb_packet_s_state_11_25),
    .I0(u_usb_device_controller_u_usb_packet_s_state[8]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[7]),
    .I2(u_usb_device_controller_u_usb_packet_s_txready),
    .I3(u_usb_device_controller_u_usb_packet_n633_44) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_11_s20 .INIT=16'h00F1;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s11  (
    .F(u_usb_device_controller_usb_transact_inst_s_sendpid_3_16),
    .I0(u_usb_device_controller_next_state[0]),
    .I1(u_usb_device_controller_next_state[2]),
    .I2(u_usb_device_controller_next_state[3]),
    .I3(u_usb_device_controller_next_state[1]) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s11 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s12  (
    .F(u_usb_device_controller_usb_transact_inst_s_sendpid_3_17),
    .I0(u_usb_device_controller_next_state[1]),
    .I1(u_usb_device_controller_next_state[2]),
    .I2(u_usb_device_controller_next_state[3]),
    .I3(u_usb_device_controller_next_state[0]) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s12 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/u_usb_packet/n640_s17  (
    .F(u_usb_device_controller_u_usb_packet_n640_22),
    .I0(u_usb_device_controller_usb_control_inst_usbc_txdat[7]),
    .I1(txdat_i_d[7]),
    .I2(txval_i_d),
    .I3(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/u_usb_packet/n640_s17 .INIT=16'hCA00;
  LUT4 \u_usb_device_controller/u_usb_packet/n640_s18  (
    .F(u_usb_device_controller_u_usb_packet_n640_23),
    .I0(u_usb_device_controller_u_usb_packet_n640_24),
    .I1(descrom_rdata_i_d[7]),
    .I2(u_usb_device_controller_u_usb_packet_n640_25),
    .I3(u_usb_device_controller_u_usb_packet_n919_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n640_s18 .INIT=16'h0700;
  LUT4 \u_usb_device_controller/u_usb_packet/n642_s17  (
    .F(u_usb_device_controller_u_usb_packet_n642_22),
    .I0(u_usb_device_controller_usb_control_inst_usbc_txdat[6]),
    .I1(txdat_i_d[6]),
    .I2(txval_i_d),
    .I3(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/u_usb_packet/n642_s17 .INIT=16'hCA00;
  LUT4 \u_usb_device_controller/u_usb_packet/n642_s18  (
    .F(u_usb_device_controller_u_usb_packet_n642_23),
    .I0(u_usb_device_controller_u_usb_packet_n640_24),
    .I1(descrom_rdata_i_d[6]),
    .I2(u_usb_device_controller_u_usb_packet_n642_24),
    .I3(u_usb_device_controller_u_usb_packet_n919_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n642_s18 .INIT=16'h0700;
  LUT4 \u_usb_device_controller/u_usb_packet/n644_s17  (
    .F(u_usb_device_controller_u_usb_packet_n644_22),
    .I0(u_usb_device_controller_u_usb_packet_n644_24),
    .I1(descrom_rdata_i_d[5]),
    .I2(u_usb_device_controller_usb_control_inst_n1649_18),
    .I3(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/u_usb_packet/n644_s17 .INIT=16'hCA00;
  LUT4 \u_usb_device_controller/u_usb_packet/n644_s18  (
    .F(u_usb_device_controller_u_usb_packet_n644_23),
    .I0(u_usb_device_controller_usb_control_inst_n2896_7),
    .I1(descrom_rdata_i_d[5]),
    .I2(u_usb_device_controller_u_usb_packet_n644_25),
    .I3(u_usb_device_controller_u_usb_packet_n919_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n644_s18 .INIT=16'h0700;
  LUT4 \u_usb_device_controller/u_usb_packet/n646_s16  (
    .F(u_usb_device_controller_u_usb_packet_n646_21),
    .I0(u_usb_device_controller_u_usb_packet_n646_24),
    .I1(descrom_rdata_i_d[4]),
    .I2(u_usb_device_controller_usb_control_inst_n1649_18),
    .I3(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/u_usb_packet/n646_s16 .INIT=16'hCA00;
  LUT3 \u_usb_device_controller/u_usb_packet/n646_s17  (
    .F(u_usb_device_controller_u_usb_packet_n646_22),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(txdat_i_d[4]),
    .I2(u_usb_device_controller_u_usb_packet_n919_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n646_s17 .INIT=8'hB0;
  LUT4 \u_usb_device_controller/u_usb_packet/n646_s18  (
    .F(u_usb_device_controller_u_usb_packet_n646_23),
    .I0(descrom_rdata_i_d[4]),
    .I1(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I2(u_usb_device_controller_u_usb_packet_n328_17),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_5_10) 
);
defparam \u_usb_device_controller/u_usb_packet/n646_s18 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/u_usb_packet/n650_s17  (
    .F(u_usb_device_controller_u_usb_packet_n650_22),
    .I0(u_usb_device_controller_u_usb_packet_n650_25),
    .I1(descrom_rdata_i_d[2]),
    .I2(u_usb_device_controller_usb_control_inst_n1649_18),
    .I3(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/u_usb_packet/n650_s17 .INIT=16'hCA00;
  LUT4 \u_usb_device_controller/u_usb_packet/n650_s18  (
    .F(u_usb_device_controller_u_usb_packet_n650_23),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(txdat_i_d[2]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[5]),
    .I3(u_usb_device_controller_usb_transact_inst_n1091_50) 
);
defparam \u_usb_device_controller/u_usb_packet/n650_s18 .INIT=16'h000B;
  LUT4 \u_usb_device_controller/u_usb_packet/n650_s19  (
    .F(u_usb_device_controller_u_usb_packet_n650_24),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(descrom_rdata_i_d[2]),
    .I2(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_5_10) 
);
defparam \u_usb_device_controller/u_usb_packet/n650_s19 .INIT=16'h7000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1672_s43  (
    .F(u_usb_device_controller_usb_control_inst_n1672_47),
    .I0(u_usb_device_controller_usbc_dsclen_1_15),
    .I1(u_usb_device_controller_usbc_dsclen_2_14),
    .I2(u_usb_device_controller_usbc_dsclen_1_14),
    .I3(u_usb_device_controller_usbc_dsclen_2_15) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s43 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/usb_control_inst/n1672_s44  (
    .F(u_usb_device_controller_usb_control_inst_n1672_48),
    .I0(u_usb_device_controller_usbc_dsclen_6_15),
    .I1(u_usb_device_controller_usbc_dsclen_4_15),
    .I2(u_usb_device_controller_usbc_dsclen_4_14),
    .I3(u_usb_device_controller_usbc_dsclen_6_14) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s44 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/usb_control_inst/n1672_s45  (
    .F(u_usb_device_controller_usb_control_inst_n1672_49),
    .I0(u_usb_device_controller_usbc_dsclen_3_14),
    .I1(u_usb_device_controller_usbc_dsclen_5_14),
    .I2(u_usb_device_controller_usbc_dsclen_7_14),
    .I3(u_usb_device_controller_usbc_dsclen_0_15) 
);
defparam \u_usb_device_controller/usb_control_inst/n1672_s45 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/usb_control_inst/n1680_s44  (
    .F(u_usb_device_controller_usb_control_inst_n1680_48),
    .I0(u_usb_device_controller_usb_control_inst_s_test_sel),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I3(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1680_s44 .INIT=16'hC07F;
  LUT2 \u_usb_device_controller/usb_control_inst/n1686_s39  (
    .F(u_usb_device_controller_usb_control_inst_n1686_43),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I1(u_usb_device_controller_usb_control_inst_s_answerlen_7_11) 
);
defparam \u_usb_device_controller/usb_control_inst/n1686_s39 .INIT=4'h4;
  LUT4 \u_usb_device_controller/usb_control_inst/n1686_s40  (
    .F(u_usb_device_controller_usb_control_inst_n1686_44),
    .I0(u_usb_device_controller_usb_control_inst_n1676_39),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I2(u_usb_device_controller_usb_control_inst_n1686_48),
    .I3(u_usb_device_controller_usb_control_inst_s_setupptr[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1686_s40 .INIT=16'h770F;
  LUT4 \u_usb_device_controller/usb_control_inst/n1690_s35  (
    .F(u_usb_device_controller_usb_control_inst_n1690_39),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]),
    .I3(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1690_s35 .INIT=16'h1E47;
  LUT4 \u_usb_device_controller/u_usb_packet/n628_s45  (
    .F(u_usb_device_controller_u_usb_packet_n628_49),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]) 
);
defparam \u_usb_device_controller/u_usb_packet/n628_s45 .INIT=16'h1428;
  LUT4 \u_usb_device_controller/u_usb_packet/n628_s46  (
    .F(u_usb_device_controller_u_usb_packet_n628_50),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]) 
);
defparam \u_usb_device_controller/u_usb_packet/n628_s46 .INIT=16'h1428;
  LUT4 \u_usb_device_controller/u_usb_packet/n633_s39  (
    .F(u_usb_device_controller_u_usb_packet_n633_43),
    .I0(u_usb_device_controller_u_usb_packet_s_state[5]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[6]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[4]),
    .I3(u_usb_device_controller_u_usb_packet_n800_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n633_s39 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/u_usb_packet/n633_s40  (
    .F(u_usb_device_controller_u_usb_packet_n633_44),
    .I0(u_usb_device_controller_u_usb_packet_s_state[0]),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I2(u_usb_device_controller_u_usb_packet_s_state[1]),
    .I3(u_usb_device_controller_u_usb_packet_n1454_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n633_s40 .INIT=16'h4000;
  LUT3 \u_usb_device_controller/usb_control_inst/n1860_s28  (
    .F(u_usb_device_controller_usb_control_inst_n1860_33),
    .I0(u_usb_device_controller_usb_control_inst_n1860_34),
    .I1(u_usb_device_controller_usb_control_inst_n645),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1860_s28 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/u_usb_init/n219_s22  (
    .F(u_usb_device_controller_u_usb_init_n219_30),
    .I0(u_usb_device_controller_u_usb_init_s_chirpcnt[0]),
    .I1(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .I2(u_usb_device_controller_u_usb_init_s_linestate[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n219_s22 .INIT=8'hE7;
  LUT3 \u_usb_device_controller/n1534_s28  (
    .F(u_usb_device_controller_n1534_35),
    .I0(u_usb_device_controller_s_endpt_txcork),
    .I1(u_usb_device_controller_s_halt_in),
    .I2(u_usb_device_controller_usb_transact_inst_s_setup_2) 
);
defparam \u_usb_device_controller/n1534_s28 .INIT=8'h0D;
  LUT4 \u_usb_device_controller/usbc_dsclen_0_s15  (
    .F(u_usb_device_controller_usbc_dsclen_0_20),
    .I0(desc_strvendor_len_i_d[0]),
    .I1(desc_strserial_len_i_d[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s15 .INIT=16'h305F;
  LUT3 \u_usb_device_controller/usbc_dsclen_0_s16  (
    .F(u_usb_device_controller_usbc_dsclen_0_21),
    .I0(desc_strproduct_len_i_d[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s16 .INIT=8'h0E;
  LUT3 \u_usb_device_controller/usbc_dsclen_0_s17  (
    .F(u_usb_device_controller_usbc_dsclen_0_22),
    .I0(desc_dev_len_i_d[0]),
    .I1(u_usb_device_controller_usbc_dsclen_0_24),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s17 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usbc_dsclen_0_s18  (
    .F(u_usb_device_controller_usbc_dsclen_0_23),
    .I0(desc_hscfg_len_i_d[0]),
    .I1(desc_fscfg_len_i_d[0]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s18 .INIT=8'hCA;
  LUT2 \u_usb_device_controller/usbc_dsclen_1_s16  (
    .F(u_usb_device_controller_usbc_dsclen_1_21),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s16 .INIT=4'h8;
  LUT4 \u_usb_device_controller/usbc_dsclen_1_s17  (
    .F(u_usb_device_controller_usbc_dsclen_1_22),
    .I0(desc_fscfg_len_i_d[1]),
    .I1(desc_hscfg_len_i_d[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I3(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s17 .INIT=16'h0C0A;
  LUT4 \u_usb_device_controller/usbc_dsclen_2_s13  (
    .F(u_usb_device_controller_usbc_dsclen_2_18),
    .I0(desc_fscfg_len_i_d[2]),
    .I1(desc_hscfg_len_i_d[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I3(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_2_s13 .INIT=16'h0305;
  LUT4 \u_usb_device_controller/usbc_dsclen_2_s14  (
    .F(u_usb_device_controller_usbc_dsclen_2_19),
    .I0(desc_strproduct_len_i_d[2]),
    .I1(desc_strserial_len_i_d[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_2_s14 .INIT=16'h3500;
  LUT4 \u_usb_device_controller/usbc_dsclen_2_s15  (
    .F(u_usb_device_controller_usbc_dsclen_2_20),
    .I0(u_usb_device_controller_usb_control_inst_n1709_17),
    .I1(desc_strvendor_len_i_d[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_2_s15 .INIT=16'h0D00;
  LUT4 \u_usb_device_controller/usbc_dsclen_3_s13  (
    .F(u_usb_device_controller_usbc_dsclen_3_18),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(desc_strproduct_len_i_d[3]),
    .I2(desc_strserial_len_i_d[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1705_16) 
);
defparam \u_usb_device_controller/usbc_dsclen_3_s13 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/usbc_dsclen_3_s14  (
    .F(u_usb_device_controller_usbc_dsclen_3_19),
    .I0(desc_fscfg_len_i_d[3]),
    .I1(desc_hscfg_len_i_d[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I3(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_3_s14 .INIT=16'h0C0A;
  LUT3 \u_usb_device_controller/usbc_dsclen_3_s15  (
    .F(u_usb_device_controller_usbc_dsclen_3_20),
    .I0(desc_hscfg_len_i_d[3]),
    .I1(desc_fscfg_len_i_d[3]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_3_s15 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/usbc_dsclen_4_s14  (
    .F(u_usb_device_controller_usbc_dsclen_4_19),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(desc_strproduct_len_i_d[4]),
    .I2(desc_strserial_len_i_d[4]),
    .I3(u_usb_device_controller_usb_control_inst_n1705_16) 
);
defparam \u_usb_device_controller/usbc_dsclen_4_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/usbc_dsclen_5_s13  (
    .F(u_usb_device_controller_usbc_dsclen_5_18),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(desc_strproduct_len_i_d[5]),
    .I2(desc_strserial_len_i_d[5]),
    .I3(u_usb_device_controller_usb_control_inst_n1705_16) 
);
defparam \u_usb_device_controller/usbc_dsclen_5_s13 .INIT=16'h0777;
  LUT3 \u_usb_device_controller/usbc_dsclen_5_s14  (
    .F(u_usb_device_controller_usbc_dsclen_5_19),
    .I0(desc_fscfg_len_i_d[5]),
    .I1(desc_hscfg_len_i_d[5]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_5_s14 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usbc_dsclen_5_s15  (
    .F(u_usb_device_controller_usbc_dsclen_5_20),
    .I0(desc_hscfg_len_i_d[5]),
    .I1(desc_fscfg_len_i_d[5]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_5_s15 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/usbc_dsclen_6_s13  (
    .F(u_usb_device_controller_usbc_dsclen_6_18),
    .I0(desc_strvendor_len_i_d[6]),
    .I1(desc_strserial_len_i_d[6]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_6_s13 .INIT=16'h305F;
  LUT3 \u_usb_device_controller/usbc_dsclen_6_s14  (
    .F(u_usb_device_controller_usbc_dsclen_6_19),
    .I0(desc_strproduct_len_i_d[6]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_6_s14 .INIT=8'h0E;
  LUT3 \u_usb_device_controller/usbc_dsclen_6_s15  (
    .F(u_usb_device_controller_usbc_dsclen_6_20),
    .I0(desc_dev_len_i_d[6]),
    .I1(u_usb_device_controller_usbc_dsclen_6_21),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_6_s15 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/usbc_dsclen_7_s13  (
    .F(u_usb_device_controller_usbc_dsclen_7_18),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(desc_strproduct_len_i_d[7]),
    .I2(desc_strserial_len_i_d[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1705_16) 
);
defparam \u_usb_device_controller/usbc_dsclen_7_s13 .INIT=16'h0777;
  LUT3 \u_usb_device_controller/usbc_dsclen_7_s14  (
    .F(u_usb_device_controller_usbc_dsclen_7_19),
    .I0(desc_fscfg_len_i_d[7]),
    .I1(desc_hscfg_len_i_d[7]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_7_s14 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/usbc_dsclen_7_s15  (
    .F(u_usb_device_controller_usbc_dsclen_7_20),
    .I0(desc_hscfg_len_i_d[7]),
    .I1(desc_fscfg_len_i_d[7]),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_7_s15 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/descrom_start_0_s14  (
    .F(u_usb_device_controller_descrom_start_0_19),
    .I0(u_usb_device_controller_descrom_start_0_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[0]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_0_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/descrom_start_1_s14  (
    .F(u_usb_device_controller_descrom_start_1_19),
    .I0(u_usb_device_controller_descrom_start_1_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[1]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_1_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/descrom_start_2_s14  (
    .F(u_usb_device_controller_descrom_start_2_19),
    .I0(u_usb_device_controller_descrom_start_2_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[2]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_2_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/descrom_start_3_s14  (
    .F(u_usb_device_controller_descrom_start_3_19),
    .I0(u_usb_device_controller_descrom_start_3_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[3]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_3_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/descrom_start_4_s14  (
    .F(u_usb_device_controller_descrom_start_4_19),
    .I0(u_usb_device_controller_descrom_start_4_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[4]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_4_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/descrom_start_5_s14  (
    .F(u_usb_device_controller_descrom_start_5_19),
    .I0(u_usb_device_controller_descrom_start_5_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[5]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_5_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/descrom_start_6_s14  (
    .F(u_usb_device_controller_descrom_start_6_19),
    .I0(u_usb_device_controller_descrom_start_6_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[6]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_6_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/descrom_start_7_s14  (
    .F(u_usb_device_controller_descrom_start_7_19),
    .I0(u_usb_device_controller_descrom_start_7_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[7]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_7_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/descrom_start_8_s14  (
    .F(u_usb_device_controller_descrom_start_8_19),
    .I0(u_usb_device_controller_descrom_start_8_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[8]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_8_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/descrom_start_9_s14  (
    .F(u_usb_device_controller_descrom_start_9_19),
    .I0(u_usb_device_controller_descrom_start_9_20),
    .I1(u_usb_device_controller_usb_control_inst_n1876_9),
    .I2(desc_strserial_addr_i_d[9]),
    .I3(u_usb_device_controller_descrom_start_0_23) 
);
defparam \u_usb_device_controller/descrom_start_9_s14 .INIT=16'h0777;
  LUT4 \u_usb_device_controller/u_usb_packet/n771_s9  (
    .F(u_usb_device_controller_u_usb_packet_n771_13),
    .I0(u_usb_device_controller_u_usb_packet_n771_15),
    .I1(descrom_rdata_i_d[3]),
    .I2(u_usb_device_controller_usb_control_inst_n1649_18),
    .I3(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s9 .INIT=16'hCA00;
  LUT4 \u_usb_device_controller/u_usb_packet/n771_s10  (
    .F(u_usb_device_controller_u_usb_packet_n771_14),
    .I0(u_usb_device_controller_usb_control_inst_n2896_7),
    .I1(descrom_rdata_i_d[3]),
    .I2(u_usb_device_controller_u_usb_packet_n771_16),
    .I3(u_usb_device_controller_u_usb_packet_n919_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s10 .INIT=16'h0700;
  LUT3 \u_usb_device_controller/u_usb_packet/n767_s5  (
    .F(u_usb_device_controller_u_usb_packet_n767_9),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid[0]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54) 
);
defparam \u_usb_device_controller/u_usb_packet/n767_s5 .INIT=8'hE0;
  LUT4 \u_usb_device_controller/u_usb_packet/n767_s6  (
    .F(u_usb_device_controller_u_usb_packet_n767_10),
    .I0(u_usb_device_controller_u_usb_packet_s_rxerror),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I2(u_usb_device_controller_usb_transact_inst_n1565_4),
    .I3(u_usb_device_controller_u_usb_packet_n912_14) 
);
defparam \u_usb_device_controller/u_usb_packet/n767_s6 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s19  (
    .F(u_usb_device_controller_u_usb_packet_n912_22),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[0]),
    .I1(u_usb_device_controller_u_usb_packet_crc16_buf[2]),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf[3]),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf[1]) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s19 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/u_usb_packet/n912_s20  (
    .F(u_usb_device_controller_u_usb_packet_n912_23),
    .I0(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I1(u_usb_device_controller_u_usb_packet_n633_43),
    .I2(u_usb_device_controller_u_usb_packet_n912_14),
    .I3(u_usb_device_controller_u_usb_packet_crc5_buf_4_11) 
);
defparam \u_usb_device_controller/u_usb_packet/n912_s20 .INIT=16'hF400;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s38  (
    .F(u_usb_device_controller_u_usb_init_n212_46),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[1]),
    .I1(u_usb_device_controller_u_usb_init_s_timer1[3]),
    .I2(u_usb_device_controller_u_usb_init_s_timer1[6]),
    .I3(u_usb_device_controller_u_usb_init_s_timer1[11]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s38 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s39  (
    .F(u_usb_device_controller_u_usb_init_n212_47),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[2]),
    .I1(u_usb_device_controller_u_usb_init_s_timer1[9]),
    .I2(u_usb_device_controller_u_usb_init_s_timer1[10]),
    .I3(u_usb_device_controller_u_usb_init_s_timer1[13]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s39 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s40  (
    .F(u_usb_device_controller_u_usb_init_n212_48),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[5]),
    .I1(u_usb_device_controller_u_usb_init_s_timer1[7]),
    .I2(u_usb_device_controller_u_usb_init_s_timer1[4]),
    .I3(u_usb_device_controller_u_usb_init_s_timer1[8]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s40 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s41  (
    .F(u_usb_device_controller_u_usb_init_n212_49),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[5]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[12]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[7]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[16]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s41 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/u_usb_init/n212_s42  (
    .F(u_usb_device_controller_u_usb_init_n212_50),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[19]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[10]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[9]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s42 .INIT=8'h40;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s43  (
    .F(u_usb_device_controller_u_usb_init_n212_51),
    .I0(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[14]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[18]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[13]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s43 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s44  (
    .F(u_usb_device_controller_u_usb_init_n212_52),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[9]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[10]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[13]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[14]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s44 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s45  (
    .F(u_usb_device_controller_u_usb_init_n212_53),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[6]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[5]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[8]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[11]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s45 .INIT=16'h0007;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s46  (
    .F(u_usb_device_controller_u_usb_init_n212_54),
    .I0(u_usb_device_controller_u_usb_init_n215_63),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[12]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[16]),
    .I3(u_usb_device_controller_u_usb_init_n212_55) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s46 .INIT=16'hD000;
  LUT3 \u_usb_device_controller/u_usb_init/n215_s54  (
    .F(u_usb_device_controller_u_usb_init_n215_61),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[15]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[17]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[6]) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s54 .INIT=8'h10;
  LUT4 \u_usb_device_controller/u_usb_init/n215_s55  (
    .F(u_usb_device_controller_u_usb_init_n215_62),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[16]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[18]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[8]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[12]) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s55 .INIT=16'h1000;
  LUT2 \u_usb_device_controller/u_usb_init/n215_s56  (
    .F(u_usb_device_controller_u_usb_init_n215_63),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[13]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[14]) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s56 .INIT=4'h1;
  LUT2 \u_usb_device_controller/u_usb_packet/n328_s21  (
    .F(u_usb_device_controller_u_usb_packet_n328_25),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(txdat_i_d[1]) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s21 .INIT=4'h4;
  LUT2 \u_usb_device_controller/u_usb_init/s_state_3_s11  (
    .F(u_usb_device_controller_u_usb_init_s_state_3_16),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[7]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[11]) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s11 .INIT=4'h4;
  LUT4 \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s11  (
    .F(u_usb_device_controller_u_usb_init_s_chirpcnt_2_15),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[4]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[5]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[12]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[16]) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s11 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/u_usb_packet/n640_s19  (
    .F(u_usb_device_controller_u_usb_packet_n640_24),
    .I0(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I1(u_usb_device_controller_usb_control_inst_s_answerptr_5_10),
    .I2(u_usb_device_controller_usb_control_inst_n1649_18),
    .I3(u_usb_device_controller_u_usb_packet_n328_17) 
);
defparam \u_usb_device_controller/u_usb_packet/n640_s19 .INIT=16'hF800;
  LUT2 \u_usb_device_controller/u_usb_packet/n640_s20  (
    .F(u_usb_device_controller_u_usb_packet_n640_25),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(txdat_i_d[7]) 
);
defparam \u_usb_device_controller/u_usb_packet/n640_s20 .INIT=4'h4;
  LUT2 \u_usb_device_controller/u_usb_packet/n642_s19  (
    .F(u_usb_device_controller_u_usb_packet_n642_24),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(txdat_i_d[6]) 
);
defparam \u_usb_device_controller/u_usb_packet/n642_s19 .INIT=4'h4;
  LUT3 \u_usb_device_controller/u_usb_packet/n644_s19  (
    .F(u_usb_device_controller_u_usb_packet_n644_24),
    .I0(u_usb_device_controller_usb_control_inst_usbc_txdat[5]),
    .I1(txdat_i_d[5]),
    .I2(txval_i_d) 
);
defparam \u_usb_device_controller/u_usb_packet/n644_s19 .INIT=8'hCA;
  LUT2 \u_usb_device_controller/u_usb_packet/n644_s20  (
    .F(u_usb_device_controller_u_usb_packet_n644_25),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(txdat_i_d[5]) 
);
defparam \u_usb_device_controller/u_usb_packet/n644_s20 .INIT=4'h4;
  LUT3 \u_usb_device_controller/u_usb_packet/n646_s19  (
    .F(u_usb_device_controller_u_usb_packet_n646_24),
    .I0(u_usb_device_controller_usb_control_inst_usbc_txdat[4]),
    .I1(txdat_i_d[4]),
    .I2(txval_i_d) 
);
defparam \u_usb_device_controller/u_usb_packet/n646_s19 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/u_usb_packet/n650_s20  (
    .F(u_usb_device_controller_u_usb_packet_n650_25),
    .I0(u_usb_device_controller_usb_control_inst_usbc_txdat[2]),
    .I1(txdat_i_d[2]),
    .I2(txval_i_d) 
);
defparam \u_usb_device_controller/u_usb_packet/n650_s20 .INIT=8'hCA;
  LUT4 \u_usb_device_controller/usb_control_inst/n1860_s29  (
    .F(u_usb_device_controller_usb_control_inst_n1860_34),
    .I0(u_usb_device_controller_halt_out[1]),
    .I1(u_usb_device_controller_halt_in[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1860_s29 .INIT=16'hCA00;
  LUT4 \u_usb_device_controller/usbc_dsclen_0_s19  (
    .F(u_usb_device_controller_usbc_dsclen_0_24),
    .I0(desc_fscfg_len_i_d[0]),
    .I1(desc_hscfg_len_i_d[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I3(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s19 .INIT=16'h0C0A;
  LUT4 \u_usb_device_controller/usbc_dsclen_6_s16  (
    .F(u_usb_device_controller_usbc_dsclen_6_21),
    .I0(desc_fscfg_len_i_d[6]),
    .I1(desc_hscfg_len_i_d[6]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I3(u_usb_device_controller_u_usb_init_highspeed_o_d) 
);
defparam \u_usb_device_controller/usbc_dsclen_6_s16 .INIT=16'h0C0A;
  LUT3 \u_usb_device_controller/descrom_start_0_s15  (
    .F(u_usb_device_controller_descrom_start_0_20),
    .I0(desc_strlang_addr_i_d[0]),
    .I1(desc_strvendor_addr_i_d[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_0_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/descrom_start_1_s15  (
    .F(u_usb_device_controller_descrom_start_1_20),
    .I0(desc_strlang_addr_i_d[1]),
    .I1(desc_strvendor_addr_i_d[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_1_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/descrom_start_2_s15  (
    .F(u_usb_device_controller_descrom_start_2_20),
    .I0(desc_strlang_addr_i_d[2]),
    .I1(desc_strvendor_addr_i_d[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_2_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/descrom_start_3_s15  (
    .F(u_usb_device_controller_descrom_start_3_20),
    .I0(desc_strlang_addr_i_d[3]),
    .I1(desc_strvendor_addr_i_d[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_3_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/descrom_start_4_s15  (
    .F(u_usb_device_controller_descrom_start_4_20),
    .I0(desc_strlang_addr_i_d[4]),
    .I1(desc_strvendor_addr_i_d[4]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_4_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/descrom_start_5_s15  (
    .F(u_usb_device_controller_descrom_start_5_20),
    .I0(desc_strlang_addr_i_d[5]),
    .I1(desc_strvendor_addr_i_d[5]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_5_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/descrom_start_6_s15  (
    .F(u_usb_device_controller_descrom_start_6_20),
    .I0(desc_strlang_addr_i_d[6]),
    .I1(desc_strvendor_addr_i_d[6]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_6_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/descrom_start_7_s15  (
    .F(u_usb_device_controller_descrom_start_7_20),
    .I0(desc_strlang_addr_i_d[7]),
    .I1(desc_strvendor_addr_i_d[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_7_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/descrom_start_8_s15  (
    .F(u_usb_device_controller_descrom_start_8_20),
    .I0(desc_strlang_addr_i_d[8]),
    .I1(desc_strvendor_addr_i_d[8]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_8_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/descrom_start_9_s15  (
    .F(u_usb_device_controller_descrom_start_9_20),
    .I0(desc_strlang_addr_i_d[9]),
    .I1(desc_strvendor_addr_i_d[9]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/descrom_start_9_s15 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/u_usb_packet/n771_s11  (
    .F(u_usb_device_controller_u_usb_packet_n771_15),
    .I0(u_usb_device_controller_usb_control_inst_usbc_txdat[3]),
    .I1(txdat_i_d[3]),
    .I2(txval_i_d) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s11 .INIT=8'hCA;
  LUT2 \u_usb_device_controller/u_usb_packet/n771_s12  (
    .F(u_usb_device_controller_u_usb_packet_n771_16),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(txdat_i_d[3]) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s12 .INIT=4'h4;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s47  (
    .F(u_usb_device_controller_u_usb_init_n212_55),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[15]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[17]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[18]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[19]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s47 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1080_s48  (
    .F(u_usb_device_controller_usb_transact_inst_n1080_53),
    .I0(u_usb_device_controller_usb_transact_inst_n1157_27),
    .I1(u_usb_device_controller_usb_transact_inst_n1041_4),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[9]),
    .I3(u_usb_device_controller_usb_transact_inst_s_state[10]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1080_s48 .INIT=16'h0008;
  LUT3 \u_usb_device_controller/n1266_s2  (
    .F(u_usb_device_controller_n1266),
    .I0(txdat_len_i_d[10]),
    .I1(txdat_len_i_d[11]),
    .I2(txdat_len_i_d[5]) 
);
defparam \u_usb_device_controller/n1266_s2 .INIT=8'h10;
  LUT4 \u_usb_device_controller/n1595_s16  (
    .F(u_usb_device_controller_n1595_23),
    .I0(u_usb_device_controller_s_bufptr[9]),
    .I1(u_usb_device_controller_n1601_23),
    .I2(u_usb_device_controller_s_bufptr[7]),
    .I3(u_usb_device_controller_s_bufptr[8]) 
);
defparam \u_usb_device_controller/n1595_s16 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/n1601_s16  (
    .F(u_usb_device_controller_n1601_23),
    .I0(u_usb_device_controller_s_bufptr[6]),
    .I1(u_usb_device_controller_n1607_23),
    .I2(u_usb_device_controller_s_bufptr[4]),
    .I3(u_usb_device_controller_s_bufptr[5]) 
);
defparam \u_usb_device_controller/n1601_s16 .INIT=16'h8000;
  LUT3 \u_usb_device_controller/usb_control_inst/n1680_s45  (
    .F(u_usb_device_controller_usb_control_inst_n1680_50),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]),
    .I2(u_usb_device_controller_n2024_7) 
);
defparam \u_usb_device_controller/usb_control_inst/n1680_s45 .INIT=8'h10;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_7_s5  (
    .F(u_usb_device_controller_utmi_dataout_o_d_7_10),
    .I0(u_usb_device_controller_utmi_dataout_o_d_7_8),
    .I1(u_usb_device_controller_usb_control_inst_usbc_testmode[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_testmode[6]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_testmode[7]) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_7_s5 .INIT=16'h0002;
  LUT4 \u_usb_device_controller/test_packet_inst/n315_s5  (
    .F(u_usb_device_controller_test_packet_inst_n315_10),
    .I0(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[2]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I3(u_usb_device_controller_test_packet_inst_test_data_val_9) 
);
defparam \u_usb_device_controller/test_packet_inst/n315_s5 .INIT=16'hEF00;
  LUT3 \u_usb_device_controller/u_usb_init/n215_s57  (
    .F(u_usb_device_controller_u_usb_init_n215_65),
    .I0(u_usb_device_controller_u_usb_init_n212_59),
    .I1(u_usb_device_controller_u_usb_init_s_state_3_12),
    .I2(u_usb_device_controller_u_usb_init_s_state_0_4) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s57 .INIT=8'h45;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s48  (
    .F(u_usb_device_controller_u_usb_init_n212_57),
    .I0(u_usb_device_controller_u_usb_init_n212_41),
    .I1(u_usb_device_controller_u_usb_init_s_timer1[0]),
    .I2(u_usb_device_controller_u_usb_init_n212_47),
    .I3(u_usb_device_controller_u_usb_init_n212_48) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s48 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s49  (
    .F(u_usb_device_controller_u_usb_init_n212_59),
    .I0(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I1(u_usb_device_controller_u_usb_init_n215_58),
    .I2(u_usb_device_controller_u_usb_init_s_chirpcnt_2_13),
    .I3(u_usb_device_controller_u_usb_init_n212_49) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s49 .INIT=16'h1555;
  LUT4 \u_usb_device_controller/u_usb_init/n215_s58  (
    .F(u_usb_device_controller_u_usb_init_n215_67),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[7]),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[13]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[14]) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s58 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/u_usb_init/n215_s59  (
    .F(u_usb_device_controller_u_usb_init_n215_69),
    .I0(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I2(u_usb_device_controller_u_usb_init_n216_53),
    .I3(u_usb_device_controller_u_usb_init_n414_4) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s59 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_3_s12  (
    .F(u_usb_device_controller_u_usb_init_s_state_3_18),
    .I0(u_usb_device_controller_u_usb_init_s_timer2[15]),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[17]),
    .I2(u_usb_device_controller_u_usb_init_s_timer2[7]),
    .I3(u_usb_device_controller_u_usb_init_s_timer2[11]) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_3_s12 .INIT=16'h0800;
  LUT3 \u_usb_device_controller/u_usb_packet/crc5_buf_4_s8  (
    .F(u_usb_device_controller_u_usb_packet_crc5_buf_4_13),
    .I0(u_usb_device_controller_u_usb_packet_s_rxerror),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I2(u_usb_device_controller_u_usb_packet_n579_20) 
);
defparam \u_usb_device_controller/u_usb_packet/crc5_buf_4_s8 .INIT=8'h40;
  LUT3 \u_usb_device_controller/u_usb_packet/n328_s22  (
    .F(u_usb_device_controller_u_usb_packet_n328_27),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(txdat_i_d[0]),
    .I2(u_usb_device_controller_u_usb_packet_n626_41) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s22 .INIT=8'hB0;
  LUT4 \u_usb_device_controller/u_usb_packet/n624_s30  (
    .F(u_usb_device_controller_u_usb_packet_n624),
    .I0(u_usb_device_controller_u_usb_packet_n328_10),
    .I1(u_usb_device_controller_u_usb_packet_n328_11),
    .I2(u_usb_device_controller_u_usb_packet_n800_6),
    .I3(u_usb_device_controller_u_usb_packet_n624_37) 
);
defparam \u_usb_device_controller/u_usb_packet/n624_s30 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/u_usb_packet/n615_s44  (
    .F(u_usb_device_controller_u_usb_packet_n615_49),
    .I0(u_usb_device_controller_u_usb_packet_n800_9),
    .I1(u_usb_device_controller_u_usb_packet_s_state[4]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[5]),
    .I3(u_usb_device_controller_u_usb_packet_s_state[6]) 
);
defparam \u_usb_device_controller/u_usb_packet/n615_s44 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/u_usb_packet/n767_s7  (
    .F(u_usb_device_controller_u_usb_packet_n767_12),
    .I0(u_usb_device_controller_u_usb_packet_n328_17),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid[0]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[9]),
    .I3(u_usb_device_controller_usb_transact_inst_n1091_54) 
);
defparam \u_usb_device_controller/u_usb_packet/n767_s7 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/u_usb_packet/n768_s2  (
    .F(u_usb_device_controller_u_usb_packet_n768),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[0]),
    .I1(u_usb_device_controller_u_usb_packet_n912_9),
    .I2(u_usb_device_controller_u_usb_packet_n767_6),
    .I3(u_usb_device_controller_u_usb_packet_n776_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n768_s2 .INIT=16'h96FF;
  LUT4 \u_usb_device_controller/u_usb_packet/n648_s13  (
    .F(u_usb_device_controller_u_usb_packet_n648),
    .I0(u_usb_device_controller_u_usb_packet_n782_5),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout[3]),
    .I2(u_usb_device_controller_u_usb_packet_n782_6),
    .I3(u_usb_device_controller_u_usb_packet_n782_7) 
);
defparam \u_usb_device_controller/u_usb_packet/n648_s13 .INIT=16'hF4FF;
  LUT4 \u_usb_device_controller/u_usb_packet/n654_s14  (
    .F(u_usb_device_controller_u_usb_packet_n654),
    .I0(u_usb_device_controller_u_usb_packet_n785_6),
    .I1(u_usb_device_controller_u_usb_packet_n328_11),
    .I2(u_usb_device_controller_u_usb_packet_n785_7),
    .I3(u_usb_device_controller_u_usb_packet_n654_18) 
);
defparam \u_usb_device_controller/u_usb_packet/n654_s14 .INIT=16'h8FFF;
  LUT3 \u_usb_device_controller/usb_control_inst/n1655_s13  (
    .F(u_usb_device_controller_usb_control_inst_n1655_18),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1655_s13 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_control_inst/s_setupptr_2_s7  (
    .F(u_usb_device_controller_usb_control_inst_s_setupptr_2_12),
    .I0(u_usb_device_controller_usb_control_inst_s_answerptr_5_10),
    .I1(u_usb_device_controller_usb_control_inst_n1670_43),
    .I2(u_usb_device_controller_usb_control_inst_s_interface_set_8),
    .I3(u_usb_device_controller_usb_control_inst_n1682_39) 
);
defparam \u_usb_device_controller/usb_control_inst/s_setupptr_2_s7 .INIT=16'hFE00;
  LUT4 \u_usb_device_controller/usb_control_inst/n1678_s41  (
    .F(u_usb_device_controller_usb_control_inst_n1678_46),
    .I0(u_usb_device_controller_usb_transact_inst_txpop_o_d_9),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerlen[0]),
    .I3(u_usb_device_controller_usb_transact_inst_txpop_o_d_5) 
);
defparam \u_usb_device_controller/usb_control_inst/n1678_s41 .INIT=16'h5400;
  LUT3 \u_usb_device_controller/usb_control_inst/n1761_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1761_16),
    .I0(u_usb_device_controller_usb_control_inst_n1876_13),
    .I1(u_usb_device_controller_usb_control_inst_s_test_sel),
    .I2(u_usb_device_controller_usb_control_inst_n2902_5) 
);
defparam \u_usb_device_controller/usb_control_inst/n1761_s11 .INIT=8'h20;
  LUT3 \u_usb_device_controller/usb_control_inst/n1709_s14  (
    .F(u_usb_device_controller_usb_control_inst_n1709_19),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1709_s14 .INIT=8'h20;
  LUT3 \u_usb_device_controller/usb_control_inst/n1909_s2  (
    .F(u_usb_device_controller_usb_control_inst_n1909),
    .I0(u_usb_device_controller_usb_control_inst_s_test_sel),
    .I1(u_usb_device_controller_usb_control_inst_n2902_5),
    .I2(u_usb_device_controller_usb_control_inst_n1876_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1909_s2 .INIT=8'h80;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1099_s44  (
    .F(u_usb_device_controller_usb_transact_inst_n1099_49),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1099_s44 .INIT=8'h20;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s13  (
    .F(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[15]),
    .I1(u_usb_device_controller_usb_transact_inst_n1124_28),
    .I2(u_usb_device_controller_usb_transact_inst_wait_count[13]),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[14]) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s13 .INIT=16'h0004;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1124_s21  (
    .F(u_usb_device_controller_usb_transact_inst_n1124_28),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[12]),
    .I1(u_usb_device_controller_usb_transact_inst_n1133_26),
    .I2(u_usb_device_controller_usb_transact_inst_wait_count[10]),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[11]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1124_s21 .INIT=16'h0004;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1138_s29  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_35),
    .I0(u_usb_device_controller_usb_transact_inst_n1146_22),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[4]),
    .I2(u_usb_device_controller_usb_transact_inst_wait_count[5]),
    .I3(u_usb_device_controller_usb_transact_inst_wait_count[6]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s29 .INIT=16'h0002;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1138_s30  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_37),
    .I0(u_usb_device_controller_usb_transact_inst_n1565_5),
    .I1(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I2(u_usb_device_controller_usb_transact_inst_n1064_16),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_24) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s30 .INIT=16'h0004;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1136_s22  (
    .F(u_usb_device_controller_usb_transact_inst_n1136_29),
    .I0(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I1(u_usb_device_controller_usb_transact_inst_n1064_16),
    .I2(u_usb_device_controller_usb_transact_inst_n1138_24) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1136_s22 .INIT=8'h01;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1138_s31  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_39),
    .I0(u_usb_device_controller_usb_transact_inst_wait_count[7]),
    .I1(u_usb_device_controller_usb_transact_inst_wait_count[8]),
    .I2(u_usb_device_controller_usb_transact_inst_n1138_35) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s31 .INIT=8'h10;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1565_s5  (
    .F(u_usb_device_controller_usb_transact_inst_n1565),
    .I0(u_usb_device_controller_usb_transact_inst_n1565_4),
    .I1(u_usb_device_controller_usb_transact_inst_n1565_5),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I3(u_usb_device_controller_usb_transact_inst_n1565_7) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1565_s5 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usbc_dsclen_0_s20  (
    .F(u_usb_device_controller_usbc_dsclen_0),
    .I0(u_usb_device_controller_usbc_dsclen_0_28),
    .I1(u_usb_device_controller_usbc_dsclen_0_18),
    .I2(u_usb_device_controller_usbc_dsclen_0_19),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s20 .INIT=16'h0511;
  LUT4 \u_usb_device_controller/usbc_dsclen_6_s17  (
    .F(u_usb_device_controller_usbc_dsclen_6),
    .I0(u_usb_device_controller_usbc_dsclen_0_28),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[2]),
    .I2(u_usb_device_controller_usbc_dsclen_6_16),
    .I3(u_usb_device_controller_usbc_dsclen_6_15) 
);
defparam \u_usb_device_controller/usbc_dsclen_6_s17 .INIT=16'h0045;
  LUT4 \u_usb_device_controller/n1607_s16  (
    .F(u_usb_device_controller_n1607_23),
    .I0(u_usb_device_controller_s_bufptr[2]),
    .I1(u_usb_device_controller_s_bufptr[3]),
    .I2(u_usb_device_controller_s_bufptr[0]),
    .I3(u_usb_device_controller_s_bufptr[1]) 
);
defparam \u_usb_device_controller/n1607_s16 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/n1611_s16  (
    .F(u_usb_device_controller_n1611),
    .I0(u_usb_device_controller_n1613_21),
    .I1(u_usb_device_controller_s_bufptr[2]),
    .I2(u_usb_device_controller_s_bufptr[0]),
    .I3(u_usb_device_controller_s_bufptr[1]) 
);
defparam \u_usb_device_controller/n1611_s16 .INIT=16'h1444;
  LUT4 \u_usb_device_controller/n1810_s3  (
    .F(u_usb_device_controller_n1810),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I3(u_usb_device_controller_s_osync) 
);
defparam \u_usb_device_controller/n1810_s3 .INIT=16'h8008;
  LUT4 \u_usb_device_controller/utmi_txvalid_o_d_s2  (
    .F(u_usb_device_controller_utmi_txvalid_o_d_6),
    .I0(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I1(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I2(u_usb_device_controller_test_packet_inst_cnt_11_12),
    .I3(u_usb_device_controller_test_packet_inst_cnt_11_13) 
);
defparam \u_usb_device_controller/utmi_txvalid_o_d_s2 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s50  (
    .F(u_usb_device_controller_u_usb_init_n212_61),
    .I0(u_usb_device_controller_u_usb_init_n212_38),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I2(u_usb_device_controller_u_usb_init_s_state[3]),
    .I3(u_usb_device_controller_u_usb_init_n212_63) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s50 .INIT=16'h00FE;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s51  (
    .F(u_usb_device_controller_u_usb_init_n212_63),
    .I0(u_usb_device_controller_u_usb_init_s_state[1]),
    .I1(u_usb_device_controller_u_usb_init_s_state[2]),
    .I2(u_usb_device_controller_u_usb_init_n215_54),
    .I3(u_usb_device_controller_u_usb_init_s_state[3]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s51 .INIT=16'hEF00;
  LUT4 \u_usb_device_controller/u_usb_init/n216_s49  (
    .F(u_usb_device_controller_u_usb_init_n216_56),
    .I0(u_usb_device_controller_u_usb_init_n215_65),
    .I1(u_usb_device_controller_u_usb_init_s_state[1]),
    .I2(u_usb_device_controller_u_usb_init_s_state[2]),
    .I3(u_usb_device_controller_u_usb_init_n216_54) 
);
defparam \u_usb_device_controller/u_usb_init/n216_s49 .INIT=16'h007F;
  LUT4 \u_usb_device_controller/u_usb_packet/n920_s5  (
    .F(u_usb_device_controller_u_usb_packet_n920_9),
    .I0(u_usb_device_controller_u_usb_init_usbp_chirpk),
    .I1(u_usb_device_controller_u_usb_packet_s_state[1]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[0]),
    .I3(u_usb_device_controller_u_usb_packet_n1454_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n920_s5 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/u_usb_packet/PHY_TXVALID_s4  (
    .F(u_usb_device_controller_u_usb_packet_PHY_TXVALID),
    .I0(u_usb_device_controller_u_usb_packet_s_state[1]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[0]),
    .I2(u_usb_device_controller_u_usb_packet_n1454_5),
    .I3(u_usb_device_controller_u_usb_packet_n919) 
);
defparam \u_usb_device_controller/u_usb_packet/PHY_TXVALID_s4 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/u_usb_packet/n1454_s3  (
    .F(u_usb_device_controller_u_usb_packet_n1454),
    .I0(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I1(u_usb_device_controller_u_usb_packet_s_state[1]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[0]),
    .I3(u_usb_device_controller_u_usb_packet_n1454_5) 
);
defparam \u_usb_device_controller/u_usb_packet/n1454_s3 .INIT=16'hBAAA;
  LUT4 \u_usb_device_controller/u_usb_packet/n620_s43  (
    .F(u_usb_device_controller_u_usb_packet_n620),
    .I0(u_usb_device_controller_u_usb_packet_s_txready),
    .I1(u_usb_device_controller_u_usb_packet_s_state[8]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[7]),
    .I3(u_usb_device_controller_u_usb_packet_s_dataout_7_9) 
);
defparam \u_usb_device_controller/u_usb_packet/n620_s43 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1091_s48  (
    .F(u_usb_device_controller_usb_transact_inst_n1091_54),
    .I0(u_usb_device_controller_u_usb_packet_s_txfirst),
    .I1(u_usb_device_controller_u_usb_packet_s_txready),
    .I2(u_usb_device_controller_u_usb_packet_n615_43),
    .I3(u_usb_device_controller_u_usb_packet_n800_9) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1091_s48 .INIT=16'hE000;
  LUT4 \u_usb_device_controller/u_usb_packet/n624_s31  (
    .F(u_usb_device_controller_u_usb_packet_n624_37),
    .I0(u_usb_device_controller_u_usb_packet_s_txfirst),
    .I1(u_usb_device_controller_u_usb_packet_s_txready),
    .I2(u_usb_device_controller_u_usb_packet_n784_20),
    .I3(u_usb_device_controller_u_usb_packet_n615_49) 
);
defparam \u_usb_device_controller/u_usb_packet/n624_s31 .INIT=16'h1F00;
  LUT3 \u_usb_device_controller/u_usb_packet/n622_s40  (
    .F(u_usb_device_controller_u_usb_packet_n622_46),
    .I0(u_usb_device_controller_u_usb_packet_s_txfirst),
    .I1(u_usb_device_controller_u_usb_packet_s_txready),
    .I2(u_usb_device_controller_u_usb_packet_n615_49) 
);
defparam \u_usb_device_controller/u_usb_packet/n622_s40 .INIT=8'hE0;
  LUT4 \u_usb_device_controller/u_usb_packet/n784_s12  (
    .F(u_usb_device_controller_u_usb_packet_n784_16),
    .I0(u_usb_device_controller_u_usb_packet_n784_20),
    .I1(u_usb_device_controller_u_usb_packet_s_dataout_7),
    .I2(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I3(u_usb_device_controller_u_usb_init_usbp_chirpk) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s12 .INIT=16'h0004;
  LUT3 \u_usb_device_controller/u_usb_packet/n626_s43  (
    .F(u_usb_device_controller_u_usb_packet_n626_48),
    .I0(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I1(u_usb_device_controller_u_usb_init_usbp_chirpk),
    .I2(u_usb_device_controller_u_usb_packet_n784_18) 
);
defparam \u_usb_device_controller/u_usb_packet/n626_s43 .INIT=8'h10;
  LUT4 \u_usb_device_controller/usb_control_inst/n1686_s43  (
    .F(u_usb_device_controller_usb_control_inst_n1686_48),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I3(u_usb_device_controller_usb_control_inst_s_answerlen_7_11) 
);
defparam \u_usb_device_controller/usb_control_inst/n1686_s43 .INIT=16'h00FE;
  LUT4 \u_usb_device_controller/usb_control_inst/s_answerlen_7_s6  (
    .F(u_usb_device_controller_usb_control_inst_s_answerlen_7_11),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerlen_7_s6 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/usb_control_inst/n2896_s5  (
    .F(u_usb_device_controller_usb_control_inst_n2896_9),
    .I0(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I1(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I2(u_usb_device_controller_u_usb_packet_n328_17),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_5_10) 
);
defparam \u_usb_device_controller/usb_control_inst/n2896_s5 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1661_s17  (
    .F(u_usb_device_controller_usb_control_inst_n1661_22),
    .I0(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[4]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[5]),
    .I3(u_usb_device_controller_usb_control_inst_n1629_4) 
);
defparam \u_usb_device_controller/usb_control_inst/n1661_s17 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/usb_control_inst/s_answerptr_5_s10  (
    .F(u_usb_device_controller_usb_control_inst_s_answerptr_5_14),
    .I0(u_usb_device_controller_usb_control_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[5]),
    .I2(u_usb_device_controller_usb_control_inst_n1629_4),
    .I3(u_usb_device_controller_usb_control_inst_n1629_5) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerptr_5_s10 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/C_CLRIN_1_s6  (
    .F(u_usb_device_controller_usb_control_inst_C_CLRIN_1_9),
    .I0(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_11),
    .I3(u_usb_device_controller_usb_control_inst_n1682_39) 
);
defparam \u_usb_device_controller/usb_control_inst/C_CLRIN_1_s6 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/s_interface_set_s7  (
    .F(u_usb_device_controller_usb_control_inst_s_interface_set),
    .I0(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I1(u_usb_device_controller_usb_control_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_7_11),
    .I3(u_usb_device_controller_usb_control_inst_s_interface_set_9) 
);
defparam \u_usb_device_controller/usb_control_inst/s_interface_set_s7 .INIT=16'hFF10;
  LUT4 \u_usb_device_controller/usb_control_inst/s_answerlen_7_s7  (
    .F(u_usb_device_controller_usb_control_inst_s_answerlen_7_13),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]) 
);
defparam \u_usb_device_controller/usb_control_inst/s_answerlen_7_s7 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1086_s43  (
    .F(u_usb_device_controller_usb_transact_inst_n1086_48),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1086_s43 .INIT=16'h0004;
  LUT3 \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s14  (
    .F(u_usb_device_controller_usb_transact_inst_s_sendpid_3_21),
    .I0(u_usb_device_controller_usb_transact_inst_s_ping),
    .I1(u_usb_device_controller_usb_transact_inst_s_in),
    .I2(u_usb_device_controller_usb_transact_inst_n1163_24) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s14 .INIT=8'hE0;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1142_s20  (
    .F(u_usb_device_controller_usb_transact_inst_n1142_25),
    .I0(u_usb_device_controller_usb_transact_inst_s_ping),
    .I1(u_usb_device_controller_usb_transact_inst_s_in),
    .I2(u_usb_device_controller_usb_transact_inst_n1074_22),
    .I3(u_usb_device_controller_usb_transact_inst_txpop_o_d_5) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1142_s20 .INIT=16'h00EF;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1148_s20  (
    .F(u_usb_device_controller_usb_transact_inst_n1148_25),
    .I0(u_usb_device_controller_usb_transact_inst_n1095_45),
    .I1(u_usb_device_controller_usb_transact_inst_n1074_22),
    .I2(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I3(u_usb_device_controller_usb_transact_inst_n1142_25) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1148_s20 .INIT=16'hF100;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1086_s44  (
    .F(u_usb_device_controller_usb_transact_inst_n1086_50),
    .I0(u_usb_device_controller_usb_transact_inst_n1072_19),
    .I1(u_usb_device_controller_usb_transact_inst_n1095_45),
    .I2(u_usb_device_controller_usb_transact_inst_n1074_22),
    .I3(u_usb_device_controller_u_usb_packet_usbp_rxact) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1086_s44 .INIT=16'hFE00;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1138_s32  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_41),
    .I0(u_usb_device_controller_usb_transact_inst_n1138_24),
    .I1(u_usb_device_controller_usb_transact_inst_n1138_25),
    .I2(u_usb_device_controller_usb_transact_inst_n1095_45),
    .I3(u_usb_device_controller_usb_transact_inst_n1074_22) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s32 .INIT=16'hFFFB;
  LUT4 \u_usb_device_controller/n1585_s2  (
    .F(u_usb_device_controller_n1585),
    .I0(u_usb_device_controller_cur_state[0]),
    .I1(u_usb_device_controller_cur_state[1]),
    .I2(u_usb_device_controller_cur_state[2]),
    .I3(u_usb_device_controller_cur_state[3]) 
);
defparam \u_usb_device_controller/n1585_s2 .INIT=16'h0008;
  LUT4 \u_usb_device_controller/n1529_s24  (
    .F(u_usb_device_controller_n1529_31),
    .I0(u_usb_device_controller_cur_state[1]),
    .I1(u_usb_device_controller_cur_state[3]),
    .I2(u_usb_device_controller_cur_state[2]),
    .I3(u_usb_device_controller_rxdat_d0_7_9) 
);
defparam \u_usb_device_controller/n1529_s24 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/rxact_o_d_s1  (
    .F(u_usb_device_controller_rxact_o_d),
    .I0(u_usb_device_controller_cur_state[0]),
    .I1(u_usb_device_controller_cur_state[1]),
    .I2(u_usb_device_controller_cur_state[3]),
    .I3(u_usb_device_controller_cur_state[2]) 
);
defparam \u_usb_device_controller/rxact_o_d_s1 .INIT=16'h0400;
  LUT4 \u_usb_device_controller/test_packet_inst/n131_s4  (
    .F(u_usb_device_controller_test_packet_inst_n131_8),
    .I0(u_usb_device_controller_test_packet_inst_cnt[5]),
    .I1(u_usb_device_controller_test_packet_inst_n133_6),
    .I2(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[4]) 
);
defparam \u_usb_device_controller/test_packet_inst/n131_s4 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/test_packet_inst/n318_s12  (
    .F(u_usb_device_controller_test_packet_inst_n318_17),
    .I0(u_usb_device_controller_test_packet_inst_cnt[3]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[0]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[1]),
    .I3(u_usb_device_controller_test_packet_inst_cnt[2]) 
);
defparam \u_usb_device_controller/test_packet_inst/n318_s12 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/u_usb_init/n210_s22  (
    .F(u_usb_device_controller_u_usb_init_n210),
    .I0(u_usb_device_controller_u_usb_init_s_state[3]),
    .I1(u_usb_device_controller_u_usb_init_s_state[2]),
    .I2(u_usb_device_controller_u_usb_init_s_state[1]),
    .I3(u_usb_device_controller_u_usb_init_s_state_0_4) 
);
defparam \u_usb_device_controller/u_usb_init/n210_s22 .INIT=16'h111F;
  LUT4 \u_usb_device_controller/u_usb_init/n209_s22  (
    .F(u_usb_device_controller_u_usb_init_n209),
    .I0(u_usb_device_controller_u_usb_init_s_state[2]),
    .I1(u_usb_device_controller_u_usb_init_s_state[3]),
    .I2(u_usb_device_controller_u_usb_init_s_state[1]),
    .I3(u_usb_device_controller_u_usb_init_s_state_0_4) 
);
defparam \u_usb_device_controller/u_usb_init/n209_s22 .INIT=16'h0009;
  LUT4 \u_usb_device_controller/u_usb_init/s_opmode_0_s3  (
    .F(u_usb_device_controller_u_usb_init_s_opmode_0),
    .I0(u_usb_device_controller_u_usb_init_s_state[2]),
    .I1(u_usb_device_controller_u_usb_init_s_state[1]),
    .I2(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I3(u_usb_device_controller_u_usb_init_s_state[3]) 
);
defparam \u_usb_device_controller/u_usb_init/s_opmode_0_s3 .INIT=16'h01FF;
  LUT3 \u_usb_device_controller/u_usb_packet/n800_s5  (
    .F(u_usb_device_controller_u_usb_packet_n800_9),
    .I0(u_usb_device_controller_u_usb_packet_s_state[2]),
    .I1(u_usb_device_controller_u_usb_packet_s_state[3]),
    .I2(u_usb_device_controller_u_usb_packet_n784_11) 
);
defparam \u_usb_device_controller/u_usb_packet/n800_s5 .INIT=8'h10;
  LUT4 \u_usb_device_controller/u_usb_packet/n784_s13  (
    .F(u_usb_device_controller_u_usb_packet_n784_18),
    .I0(u_usb_device_controller_u_usb_packet_n784_9),
    .I1(u_usb_device_controller_u_usb_packet_s_state[2]),
    .I2(u_usb_device_controller_u_usb_packet_s_state[3]),
    .I3(u_usb_device_controller_u_usb_packet_n784_11) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s13 .INIT=16'h0200;
  LUT3 \u_usb_device_controller/usb_control_inst/n1649_s18  (
    .F(u_usb_device_controller_usb_control_inst_n1649_23),
    .I0(u_usb_device_controller_usb_control_inst_n1680_50),
    .I1(u_usb_device_controller_usb_control_inst_n1474_3),
    .I2(u_usb_device_controller_usb_control_inst_n1483_3) 
);
defparam \u_usb_device_controller/usb_control_inst/n1649_s18 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1674_s37  (
    .F(u_usb_device_controller_usb_control_inst_n1674),
    .I0(u_usb_device_controller_usb_control_inst_n1672_42),
    .I1(u_usb_device_controller_usb_control_inst_n1474_3),
    .I2(u_usb_device_controller_usb_control_inst_n1483_3),
    .I3(u_usb_device_controller_usb_control_inst_n1674_39) 
);
defparam \u_usb_device_controller/usb_control_inst/n1674_s37 .INIT=16'hFF80;
  LUT3 \u_usb_device_controller/descrom_start_0_s17  (
    .F(u_usb_device_controller_descrom_start_0_23),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I1(u_usb_device_controller_usb_control_inst_n1836_11),
    .I2(u_usb_device_controller_usb_control_inst_n1705_16) 
);
defparam \u_usb_device_controller/descrom_start_0_s17 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1876_s5  (
    .F(u_usb_device_controller_usb_control_inst_n1876_9),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1836_11) 
);
defparam \u_usb_device_controller/usb_control_inst/n1876_s5 .INIT=16'h0100;
  LUT3 \u_usb_device_controller/usb_control_inst/n1836_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1836_13),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I1(u_usb_device_controller_usb_control_inst_n1836_11),
    .I2(u_usb_device_controller_usb_control_inst_n1703_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1836_s9 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1686_s44  (
    .F(u_usb_device_controller_usb_control_inst_n1686_50),
    .I0(u_usb_device_controller_usb_control_inst_n1836_8),
    .I1(u_usb_device_controller_usb_control_inst_n1836_13),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I3(u_usb_device_controller_usb_control_inst_s_setupptr[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1686_s44 .INIT=16'h0DDD;
  LUT4 \u_usb_device_controller/usb_control_inst/n1693_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1693),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[1]),
    .I3(u_usb_device_controller_usb_control_inst_n1836_15) 
);
defparam \u_usb_device_controller/usb_control_inst/n1693_s9 .INIT=16'h6A00;
  LUT4 \u_usb_device_controller/usb_control_inst/n2067_s5  (
    .F(u_usb_device_controller_usb_control_inst_n2067),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[2]),
    .I1(u_usb_device_controller_usb_control_inst_n2067_6),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I3(u_usb_device_controller_usb_control_inst_s_setupptr[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n2067_s5 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1088_s43  (
    .F(u_usb_device_controller_usb_transact_inst_n1088_48),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1088_s43 .INIT=16'h4144;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1070_s13  (
    .F(u_usb_device_controller_usb_transact_inst_n1070_18),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1070_s13 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1111_s15  (
    .F(u_usb_device_controller_usb_transact_inst_n1111),
    .I0(u_usb_device_controller_usb_transact_inst_n1064_27),
    .I1(u_usb_device_controller_usb_transact_inst_n1111_22),
    .I2(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1111_s15 .INIT=16'h0800;
  LUT4 \u_usb_device_controller/usb_transact_inst/T_PING_s3  (
    .F(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I0(u_usb_device_controller_usb_transact_inst_txpop_o_d_5),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I2(u_usb_device_controller_usb_transact_inst_n1064_16),
    .I3(u_usb_device_controller_usb_transact_inst_n1080_46) 
);
defparam \u_usb_device_controller/usb_transact_inst/T_PING_s3 .INIT=16'h0100;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1041_s4  (
    .F(u_usb_device_controller_usb_transact_inst_n1041_8),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[9]),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_28) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1041_s4 .INIT=8'h10;
  LUT4 \u_usb_device_controller/u_usb_packet/n770_s5  (
    .F(u_usb_device_controller_u_usb_packet_n770_10),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_u_usb_packet_n626_42),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54),
    .I3(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]) 
);
defparam \u_usb_device_controller/u_usb_packet/n770_s5 .INIT=16'h2F00;
  LUT4 \u_usb_device_controller/u_usb_packet/n770_s6  (
    .F(u_usb_device_controller_u_usb_packet_n770_12),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_u_usb_packet_n626_42),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54),
    .I3(u_usb_device_controller_u_usb_packet_n650_21) 
);
defparam \u_usb_device_controller/u_usb_packet/n770_s6 .INIT=16'hD000;
  LUT4 \u_usb_device_controller/u_usb_packet/n640_s21  (
    .F(u_usb_device_controller_u_usb_packet_n640_27),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_u_usb_packet_n626_42),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54),
    .I3(u_usb_device_controller_u_usb_packet_n626) 
);
defparam \u_usb_device_controller/u_usb_packet/n640_s21 .INIT=16'h002F;
  LUT4 \u_usb_device_controller/usb_transact_inst/txpop_o_d_s4  (
    .F(u_usb_device_controller_usb_transact_inst_txpop_o_d_9),
    .I0(u_usb_device_controller_u_usb_packet_n626_41),
    .I1(u_usb_device_controller_u_usb_packet_n626_42),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54),
    .I3(u_usb_device_controller_u_usb_packet_n800_6) 
);
defparam \u_usb_device_controller/usb_transact_inst/txpop_o_d_s4 .INIT=16'h002F;
  LUT3 \u_usb_device_controller/u_usb_init/s_state_2_s12  (
    .F(u_usb_device_controller_u_usb_init_s_state_2_18),
    .I0(u_usb_device_controller_u_usb_init_n212_29),
    .I1(u_usb_device_controller_u_usb_init_s_state[3]),
    .I2(u_usb_device_controller_u_usb_init_s_state[2]) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_2_s12 .INIT=8'h10;
  LUT4 \u_usb_device_controller/u_usb_init/n223_s20  (
    .F(u_usb_device_controller_u_usb_init_n223),
    .I0(u_usb_device_controller_u_usb_init_s_state[1]),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I2(u_usb_device_controller_u_usb_init_s_state[3]),
    .I3(u_usb_device_controller_u_usb_init_s_state[2]) 
);
defparam \u_usb_device_controller/u_usb_init/n223_s20 .INIT=16'h0400;
  LUT4 \u_usb_device_controller/u_usb_init/n214_s23  (
    .F(u_usb_device_controller_u_usb_init_n214),
    .I0(u_usb_device_controller_u_usb_init_s_state[1]),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I2(u_usb_device_controller_u_usb_init_s_state[3]),
    .I3(u_usb_device_controller_u_usb_init_s_state[2]) 
);
defparam \u_usb_device_controller/u_usb_init/n214_s23 .INIT=16'h0800;
  LUT4 \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s12  (
    .F(u_usb_device_controller_u_usb_init_s_chirpcnt_2),
    .I0(reset_i_d),
    .I1(u_usb_device_controller_u_usb_init_s_chirpcnt_2_8),
    .I2(u_usb_device_controller_u_usb_init_s_state[3]),
    .I3(u_usb_device_controller_u_usb_init_s_state[2]) 
);
defparam \u_usb_device_controller/u_usb_init/s_chirpcnt_2_s12 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_2_s13  (
    .F(u_usb_device_controller_u_usb_init_s_state_2_20),
    .I0(u_usb_device_controller_u_usb_init_n212_45),
    .I1(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .I2(u_usb_device_controller_u_usb_init_s_linestate[1]),
    .I3(u_usb_device_controller_u_usb_init_s_state_0_4) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_2_s13 .INIT=16'hFCAA;
  LUT4 \u_usb_device_controller/u_usb_init/n212_s52  (
    .F(u_usb_device_controller_u_usb_init_n212_65),
    .I0(u_usb_device_controller_u_usb_init_s_usb_test_en[0]),
    .I1(u_usb_device_controller_u_usb_init_s_state[1]),
    .I2(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .I3(u_usb_device_controller_u_usb_init_s_linestate[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n212_s52 .INIT=16'h0004;
  LUT4 \u_usb_device_controller/u_usb_init/n215_s60  (
    .F(u_usb_device_controller_u_usb_init_n215_71),
    .I0(u_usb_device_controller_u_usb_init_s_state[1]),
    .I1(u_usb_device_controller_u_usb_init_s_linestate[0]),
    .I2(u_usb_device_controller_u_usb_init_s_linestate[1]),
    .I3(u_usb_device_controller_u_usb_init_n215_54) 
);
defparam \u_usb_device_controller/u_usb_init/n215_s60 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/u_usb_init/s_highspeed_s6  (
    .F(u_usb_device_controller_u_usb_init_s_highspeed),
    .I0(u_usb_device_controller_u_usb_init_s_state[3]),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I2(u_usb_device_controller_u_usb_init_s_state[2]),
    .I3(u_usb_device_controller_u_usb_init_s_state[1]) 
);
defparam \u_usb_device_controller/u_usb_init/s_highspeed_s6 .INIT=16'h4144;
  LUT4 \u_usb_device_controller/u_usb_init/n414_s2  (
    .F(u_usb_device_controller_u_usb_init_n414),
    .I0(u_usb_device_controller_u_usb_init_s_state[3]),
    .I1(u_usb_device_controller_u_usb_init_s_state_0_4),
    .I2(u_usb_device_controller_u_usb_init_s_state[2]),
    .I3(u_usb_device_controller_u_usb_init_s_state[1]) 
);
defparam \u_usb_device_controller/u_usb_init/n414_s2 .INIT=16'h0400;
  LUT4 \u_usb_device_controller/u_usb_packet/crc16_buf_15_s6  (
    .F(u_usb_device_controller_u_usb_packet_crc16_buf_15_12),
    .I0(u_usb_device_controller_u_usb_packet_n919_5),
    .I1(u_usb_device_controller_u_usb_packet_n626_42),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_54),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf_15_14) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_15_s6 .INIT=16'h002F;
  LUT3 \u_usb_device_controller/usb_control_inst/n1701_s16  (
    .F(u_usb_device_controller_usb_control_inst_n1701_21),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1701_s16 .INIT=8'h02;
  LUT4 \u_usb_device_controller/usb_control_inst/n1876_s6  (
    .F(u_usb_device_controller_usb_control_inst_n1876_11),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I3(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1876_s6 .INIT=16'h0008;
  LUT4 \u_usb_device_controller/usb_control_inst/n1864_s4  (
    .F(u_usb_device_controller_usb_control_inst_n1864_8),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I1(u_usb_device_controller_usb_control_inst_s_ctlrequest[3]),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlrequest[1]),
    .I3(u_usb_device_controller_usb_control_inst_s_ctlrequest[2]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1864_s4 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/usb_control_inst/n1670_s40  (
    .F(u_usb_device_controller_usb_control_inst_n1670_45),
    .I0(u_usb_device_controller_usb_control_inst_n1649_18),
    .I1(u_usb_device_controller_usb_control_inst_s_state[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[1]),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_7_15) 
);
defparam \u_usb_device_controller/usb_control_inst/n1670_s40 .INIT=16'h4555;
  LUT4 \u_usb_device_controller/usb_control_inst/n1836_s10  (
    .F(u_usb_device_controller_usb_control_inst_n1836_15),
    .I0(u_usb_device_controller_n2393_9),
    .I1(u_usb_device_controller_usb_control_inst_s_state[0]),
    .I2(u_usb_device_controller_usb_control_inst_s_state[1]),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_7_15) 
);
defparam \u_usb_device_controller/usb_control_inst/n1836_s10 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1080_s49  (
    .F(u_usb_device_controller_usb_transact_inst_n1080_55),
    .I0(u_usb_device_controller_usb_transact_inst_n1041_4),
    .I1(u_usb_device_controller_usb_transact_inst_n1041_8),
    .I2(u_usb_device_controller_usb_transact_inst_n1041_6),
    .I3(u_usb_device_controller_usb_transact_inst_s_endpt_0_7) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1080_s49 .INIT=16'h007F;
  LUT3 \u_usb_device_controller/u_usb_packet/s_state_11_s21  (
    .F(u_usb_device_controller_u_usb_packet_s_state_11_27),
    .I0(u_usb_device_controller_u_usb_packet_s_rxerror),
    .I1(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I2(u_usb_device_controller_u_usb_packet_usbp_rxact) 
);
defparam \u_usb_device_controller/u_usb_packet/s_state_11_s21 .INIT=8'h10;
  LUT4 \u_usb_device_controller/n1240_s2  (
    .F(u_usb_device_controller_n1240),
    .I0(txcork_i_d),
    .I1(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_test_en),
    .I3(u_usb_device_controller_utmi_dataout_o_d_0_4) 
);
defparam \u_usb_device_controller/n1240_s2 .INIT=16'hEAAA;
  LUT4 \u_usb_device_controller/n503_s5  (
    .F(u_usb_device_controller_n503_10),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[3]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n503_s5 .INIT=16'h0009;
  LUT4 \u_usb_device_controller/n443_s5  (
    .F(u_usb_device_controller_n443_10),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[2]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n443_s5 .INIT=16'h0009;
  LUT4 \u_usb_device_controller/n385_s5  (
    .F(u_usb_device_controller_n385_10),
    .I0(u_usb_device_controller_osync[1]),
    .I1(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n385_s5 .INIT=16'h0009;
  LUT4 \u_usb_device_controller/isync_3_s5  (
    .F(u_usb_device_controller_isync_3),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_3_9),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_3_s5 .INIT=16'hFF10;
  LUT4 \u_usb_device_controller/isync_2_s5  (
    .F(u_usb_device_controller_isync_2),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_2_9),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_2_s5 .INIT=16'hFF10;
  LUT4 \u_usb_device_controller/isync_1_s6  (
    .F(u_usb_device_controller_isync_1),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_1_10),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_1_s6 .INIT=16'hFF10;
  LUT4 \u_usb_device_controller/n1524_s20  (
    .F(u_usb_device_controller_n1524_27),
    .I0(u_usb_device_controller_cur_state[1]),
    .I1(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I2(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I3(u_usb_device_controller_n1529_24) 
);
defparam \u_usb_device_controller/n1524_s20 .INIT=16'hAADF;
  LUT3 \u_usb_device_controller/n1534_s29  (
    .F(u_usb_device_controller_n1534_37),
    .I0(u_usb_device_controller_usb_transact_inst_T_PING_7),
    .I1(u_usb_device_controller_usb_transact_inst_s_in_valid),
    .I2(u_usb_device_controller_n1534_31) 
);
defparam \u_usb_device_controller/n1534_s29 .INIT=8'h40;
  LUT4 \u_usb_device_controller/n384_s5  (
    .F(u_usb_device_controller_n384_10),
    .I0(u_usb_device_controller_cur_state[0]),
    .I1(u_usb_device_controller_cur_state[1]),
    .I2(u_usb_device_controller_cur_state[2]),
    .I3(u_usb_device_controller_cur_state[3]) 
);
defparam \u_usb_device_controller/n384_s5 .INIT=16'h0001;
  LUT4 \u_usb_device_controller/n1519_s22  (
    .F(u_usb_device_controller_n1519_32),
    .I0(u_usb_device_controller_cur_state[2]),
    .I1(u_usb_device_controller_usb_transact_inst_s_setup_2),
    .I2(u_usb_device_controller_cur_state[0]),
    .I3(u_usb_device_controller_cur_state[1]) 
);
defparam \u_usb_device_controller/n1519_s22 .INIT=16'h0004;
  LUT4 \u_usb_device_controller/n1520_s20  (
    .F(u_usb_device_controller_n1520),
    .I0(u_usb_device_controller_cur_state[2]),
    .I1(u_usb_device_controller_cur_state[0]),
    .I2(u_usb_device_controller_cur_state[1]),
    .I3(u_usb_device_controller_cur_state[3]) 
);
defparam \u_usb_device_controller/n1520_s20 .INIT=16'h01FF;
  LUT4 \u_usb_device_controller/n1593_s16  (
    .F(u_usb_device_controller_n1593_24),
    .I0(u_usb_device_controller_cur_state[3]),
    .I1(u_usb_device_controller_cur_state[0]),
    .I2(u_usb_device_controller_cur_state[1]),
    .I3(u_usb_device_controller_n1585) 
);
defparam \u_usb_device_controller/n1593_s16 .INIT=16'hFF01;
  LUT4 \u_usb_device_controller/setup_o_d_s1  (
    .F(u_usb_device_controller_setup_o_d),
    .I0(u_usb_device_controller_cur_state[2]),
    .I1(u_usb_device_controller_cur_state[3]),
    .I2(u_usb_device_controller_cur_state[0]),
    .I3(u_usb_device_controller_cur_state[1]) 
);
defparam \u_usb_device_controller/setup_o_d_s1 .INIT=16'h0004;
  LUT3 \u_usb_device_controller/test_packet_inst/n378_s4  (
    .F(u_usb_device_controller_test_packet_inst_n378_8),
    .I0(u_usb_device_controller_test_packet_inst_test_data_6_9),
    .I1(u_usb_device_controller_test_packet_inst_cnt[4]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[5]) 
);
defparam \u_usb_device_controller/test_packet_inst/n378_s4 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1876_s7  (
    .F(u_usb_device_controller_usb_control_inst_n1876_13),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_fin),
    .I1(u_usb_device_controller_usb_control_inst_n1629_4),
    .I2(u_usb_device_controller_usb_control_inst_n1629_5),
    .I3(u_usb_device_controller_usb_control_inst_n1629_6) 
);
defparam \u_usb_device_controller/usb_control_inst/n1876_s7 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1805_s10  (
    .F(u_usb_device_controller_usb_control_inst_n1805),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_n1805_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1805_s10 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/usb_control_inst/n1775_s10  (
    .F(u_usb_device_controller_usb_control_inst_n1775),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_n1775_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1775_s10 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/test_packet_inst/n312_s8  (
    .F(u_usb_device_controller_test_packet_inst_n312_13),
    .I0(u_usb_device_controller_test_packet_inst_cnt[5]),
    .I1(u_usb_device_controller_test_packet_inst_cnt[6]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[7]),
    .I3(u_usb_device_controller_test_packet_inst_n318_13) 
);
defparam \u_usb_device_controller/test_packet_inst/n312_s8 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/test_packet_inst/test_data_val_s5  (
    .F(u_usb_device_controller_test_packet_inst_test_data_val_9),
    .I0(u_usb_device_controller_test_packet_inst_n378_8),
    .I1(u_usb_device_controller_test_packet_inst_cnt[6]),
    .I2(u_usb_device_controller_test_packet_inst_cnt[7]),
    .I3(u_usb_device_controller_test_packet_inst_n318_13) 
);
defparam \u_usb_device_controller/test_packet_inst/test_data_val_s5 .INIT=16'h0100;
  LUT4 \u_usb_device_controller/usb_control_inst/n1773_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1773),
    .I0(u_usb_device_controller_usb_control_inst_n1713_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1773_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1771_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1771),
    .I0(u_usb_device_controller_usb_control_inst_n1711_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1771_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1769_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1769),
    .I0(u_usb_device_controller_usb_control_inst_n1709_19),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1769_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1767_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1767),
    .I0(u_usb_device_controller_usb_control_inst_n1707_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1767_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1765_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1765),
    .I0(u_usb_device_controller_usb_control_inst_n1705_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1765_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1763_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1763),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1763_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1761_s12  (
    .F(u_usb_device_controller_usb_control_inst_n1761),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1761_s12 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1803_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1803),
    .I0(u_usb_device_controller_usb_control_inst_n1713_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1803_s9 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/usb_control_inst/n1801_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1801),
    .I0(u_usb_device_controller_usb_control_inst_n1711_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1801_s9 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/usb_control_inst/n1799_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1799),
    .I0(u_usb_device_controller_usb_control_inst_n1709_19),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1799_s9 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/usb_control_inst/n1797_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1797),
    .I0(u_usb_device_controller_usb_control_inst_n1707_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1797_s9 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/usb_control_inst/n1795_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1795),
    .I0(u_usb_device_controller_usb_control_inst_n1705_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1795_s9 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/usb_control_inst/n1793_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1793),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1793_s9 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/usb_control_inst/n1791_s10  (
    .F(u_usb_device_controller_usb_control_inst_n1791),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1791_s10 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/usb_control_inst/n2902_s4  (
    .F(u_usb_device_controller_usb_control_inst_n2902),
    .I0(u_usb_device_controller_usb_transact_inst_s_setup_2),
    .I1(u_usb_device_controller_usb_control_inst_n2896_9),
    .I2(u_usb_device_controller_usb_control_inst_s_test_sel),
    .I3(u_usb_device_controller_usb_control_inst_n2902_5) 
);
defparam \u_usb_device_controller/usb_control_inst/n2902_s4 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1388_s6  (
    .F(u_usb_device_controller_usb_control_inst_n1388_12),
    .I0(u_usb_device_controller_usb_control_inst_s_ctlrequest[0]),
    .I1(u_usb_device_controller_usb_transact_inst_s_setup_2),
    .I2(u_usb_device_controller_usb_control_inst_n2896_9),
    .I3(u_usb_device_controller_usb_control_inst_n1837_6) 
);
defparam \u_usb_device_controller/usb_control_inst/n1388_s6 .INIT=16'h1000;
  LUT3 \u_usb_device_controller/usb_control_inst/n1676_s36  (
    .F(u_usb_device_controller_usb_control_inst_n1676),
    .I0(u_usb_device_controller_usb_transact_inst_s_setup_2),
    .I1(u_usb_device_controller_usb_control_inst_n2896_9),
    .I2(u_usb_device_controller_usb_control_inst_n1676_39) 
);
defparam \u_usb_device_controller/usb_control_inst/n1676_s36 .INIT=8'h40;
  LUT4 \u_usb_device_controller/n1231_s4  (
    .F(u_usb_device_controller_n1231_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[15]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n1231_s4 .INIT=16'h9000;
  LUT4 \u_usb_device_controller/n1167_s4  (
    .F(u_usb_device_controller_n1167_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[14]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n1167_s4 .INIT=16'h9000;
  LUT4 \u_usb_device_controller/n1105_s4  (
    .F(u_usb_device_controller_n1105_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[13]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n1105_s4 .INIT=16'h9000;
  LUT4 \u_usb_device_controller/n1043_s4  (
    .F(u_usb_device_controller_n1043_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[12]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n1043_s4 .INIT=16'h9000;
  LUT4 \u_usb_device_controller/isync_15_s4  (
    .F(u_usb_device_controller_isync_15),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_3_9),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_15_s4 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/isync_14_s4  (
    .F(u_usb_device_controller_isync_14),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_2_9),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_14_s4 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/isync_13_s4  (
    .F(u_usb_device_controller_isync_13),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_1_10),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_13_s4 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/isync_12_s5  (
    .F(u_usb_device_controller_isync_12),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_4_10),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_12_s5 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/n743_s4  (
    .F(u_usb_device_controller_n743_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[7]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
defparam \u_usb_device_controller/n743_s4 .INIT=16'h0900;
  LUT4 \u_usb_device_controller/n681_s4  (
    .F(u_usb_device_controller_n681_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[6]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
defparam \u_usb_device_controller/n681_s4 .INIT=16'h0900;
  LUT4 \u_usb_device_controller/n621_s4  (
    .F(u_usb_device_controller_n621_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[5]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
defparam \u_usb_device_controller/n621_s4 .INIT=16'h0900;
  LUT4 \u_usb_device_controller/n561_s5  (
    .F(u_usb_device_controller_n561_10),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[4]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]) 
);
defparam \u_usb_device_controller/n561_s5 .INIT=16'h0900;
  LUT4 \u_usb_device_controller/isync_7_s4  (
    .F(u_usb_device_controller_isync_7),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I2(u_usb_device_controller_isync_3_9),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_7_s4 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/isync_6_s4  (
    .F(u_usb_device_controller_isync_6),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I2(u_usb_device_controller_isync_2_9),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_6_s4 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/isync_5_s4  (
    .F(u_usb_device_controller_isync_5),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I2(u_usb_device_controller_isync_1_10),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_5_s4 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/isync_4_s6  (
    .F(u_usb_device_controller_isync_4),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I2(u_usb_device_controller_isync_4_10),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_4_s6 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/n983_s4  (
    .F(u_usb_device_controller_n983_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[11]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n983_s4 .INIT=16'h0900;
  LUT4 \u_usb_device_controller/n921_s4  (
    .F(u_usb_device_controller_n921_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[10]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n921_s4 .INIT=16'h0900;
  LUT4 \u_usb_device_controller/n861_s4  (
    .F(u_usb_device_controller_n861_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[9]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n861_s4 .INIT=16'h0900;
  LUT4 \u_usb_device_controller/n801_s4  (
    .F(u_usb_device_controller_n801_9),
    .I0(u_usb_device_controller_usb_transact_inst_usbt_osync),
    .I1(u_usb_device_controller_osync[8]),
    .I2(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I3(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]) 
);
defparam \u_usb_device_controller/n801_s4 .INIT=16'h0900;
  LUT4 \u_usb_device_controller/isync_11_s4  (
    .F(u_usb_device_controller_isync_11),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_3_9),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_11_s4 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/isync_10_s4  (
    .F(u_usb_device_controller_isync_10),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_2_9),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_10_s4 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/isync_9_s4  (
    .F(u_usb_device_controller_isync_9),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_1_10),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_9_s4 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/isync_8_s5  (
    .F(u_usb_device_controller_isync_8),
    .I0(u_usb_device_controller_usb_transact_inst_endpt_o_d[2]),
    .I1(u_usb_device_controller_usb_transact_inst_endpt_o_d[3]),
    .I2(u_usb_device_controller_isync_4_10),
    .I3(u_usb_device_controller_n384_10) 
);
defparam \u_usb_device_controller/isync_8_s5 .INIT=16'hFF40;
  LUT4 \u_usb_device_controller/usb_control_inst/n1813_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1813),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_n1805_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1813_s9 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1783_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1783),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_n1775_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1783_s9 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1817_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1817),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_n1805_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1817_s9 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1787_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1787),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_n1775_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1787_s9 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1819_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1819),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_n1805_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1819_s9 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1789_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1789),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_n1775_13) 
);
defparam \u_usb_device_controller/usb_control_inst/n1789_s9 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1785_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1785),
    .I0(u_usb_device_controller_usb_control_inst_n1709_19),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1785_s9 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1781_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1781),
    .I0(u_usb_device_controller_usb_control_inst_n1705_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1781_s9 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1779_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1779),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1779_s9 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1777_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1777),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1777_s9 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1815_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1815),
    .I0(u_usb_device_controller_usb_control_inst_n1709_19),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1815_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1811_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1811),
    .I0(u_usb_device_controller_usb_control_inst_n1705_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1811_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1809_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1809),
    .I0(u_usb_device_controller_usb_control_inst_n1703_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1809_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1807_s9  (
    .F(u_usb_device_controller_usb_control_inst_n1807),
    .I0(u_usb_device_controller_usb_control_inst_n1701_16),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I3(u_usb_device_controller_usb_control_inst_n1761_16) 
);
defparam \u_usb_device_controller/usb_control_inst/n1807_s9 .INIT=16'h2000;
  LUT4 \u_usb_device_controller/utmi_txvalid_o_d_s3  (
    .F(u_usb_device_controller_utmi_txvalid_o_d_8),
    .I0(u_usb_device_controller_utmi_dataout_o_d_7_7),
    .I1(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I2(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I3(u_usb_device_controller_utmi_dataout_o_d_7_10) 
);
defparam \u_usb_device_controller/utmi_txvalid_o_d_s3 .INIT=16'h1555;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_1_s1  (
    .F(u_usb_device_controller_utmi_dataout_o_d[1]),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_10),
    .I3(u_usb_device_controller_utmi_dataout_o_d_1) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_1_s1 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_2_s1  (
    .F(u_usb_device_controller_utmi_dataout_o_d[2]),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_10),
    .I3(u_usb_device_controller_utmi_dataout_o_d_2) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_2_s1 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_3_s1  (
    .F(u_usb_device_controller_utmi_dataout_o_d[3]),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_10),
    .I3(u_usb_device_controller_utmi_dataout_o_d_3) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_3_s1 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_4_s1  (
    .F(u_usb_device_controller_utmi_dataout_o_d[4]),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_10),
    .I3(u_usb_device_controller_utmi_dataout_o_d_4) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_4_s1 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_5_s1  (
    .F(u_usb_device_controller_utmi_dataout_o_d[5]),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_10),
    .I3(u_usb_device_controller_utmi_dataout_o_d_5) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_5_s1 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_6_s1  (
    .F(u_usb_device_controller_utmi_dataout_o_d[6]),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_10),
    .I3(u_usb_device_controller_utmi_dataout_o_d_6) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_6_s1 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/utmi_dataout_o_d_7_s6  (
    .F(u_usb_device_controller_utmi_dataout_o_d[7]),
    .I0(u_usb_device_controller_usb_control_inst_usbc_testmode[0]),
    .I1(u_usb_device_controller_test_packet_inst_test_en_dly_Z),
    .I2(u_usb_device_controller_utmi_dataout_o_d_7_10),
    .I3(u_usb_device_controller_utmi_dataout_o_d_7) 
);
defparam \u_usb_device_controller/utmi_dataout_o_d_7_s6 .INIT=16'hFF80;
  LUT4 \u_usb_device_controller/usb_control_inst/n1652_s17  (
    .F(u_usb_device_controller_usb_control_inst_n1652_22),
    .I0(u_usb_device_controller_usb_control_inst_n1661_17),
    .I1(u_usb_device_controller_usb_control_inst_n1649_23),
    .I2(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I3(u_usb_device_controller_usb_control_inst_s_answerptr_5_14) 
);
defparam \u_usb_device_controller/usb_control_inst/n1652_s17 .INIT=16'h0777;
  LUT3 \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s14  (
    .F(u_usb_device_controller_usb_control_inst_s_sendbyte_7_19),
    .I0(u_usb_device_controller_usb_control_inst_s_sendbyte_7_15),
    .I1(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_5_14) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s14 .INIT=8'h40;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1101_s43  (
    .F(u_usb_device_controller_usb_transact_inst_n1101_48),
    .I0(u_usb_device_controller_usb_transact_inst_n1090_46),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1101_s43 .INIT=8'h40;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1070_s14  (
    .F(u_usb_device_controller_usb_transact_inst_n1070_20),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I2(u_usb_device_controller_usb_transact_inst_n1068_18) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1070_s14 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1076_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1076_24),
    .I0(u_usb_device_controller_usb_transact_inst_n1068_18),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I3(u_usb_device_controller_usb_transact_inst_s_out_valid) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1076_s17 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1163_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1163_24),
    .I0(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I1(u_usb_device_controller_usb_transact_inst_s_prevrxact),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I3(u_usb_device_controller_usb_transact_inst_n1157_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1163_s19 .INIT=16'h1000;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1068_s10  (
    .F(u_usb_device_controller_usb_transact_inst_n1068_16),
    .I0(u_usb_device_controller_usb_transact_inst_n1068_18),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I3(u_usb_device_controller_usb_transact_inst_n1064_16) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1068_s10 .INIT=16'h00BF;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1076_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1076_26),
    .I0(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I1(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I2(u_usb_device_controller_usb_transact_inst_n1074_22),
    .I3(u_usb_device_controller_usb_transact_inst_n1064_27) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1076_s18 .INIT=16'hFFF8;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1064_s17  (
    .F(u_usb_device_controller_usb_transact_inst_n1064_23),
    .I0(u_usb_device_controller_usb_transact_inst_n1064_16),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I3(u_usb_device_controller_usb_transact_inst_n1064_27) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1064_s17 .INIT=16'hFFEA;
  LUT3 \u_usb_device_controller/rxval_o_d_s0  (
    .F(u_usb_device_controller_rxval_o_d),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_rxval_d2) 
);
defparam \u_usb_device_controller/rxval_o_d_s0 .INIT=8'hE0;
  LUT3 \u_usb_device_controller/rxdat_o_d_0_s0  (
    .F(u_usb_device_controller_rxdat_o_d[0]),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_rxdat_d2[0]) 
);
defparam \u_usb_device_controller/rxdat_o_d_0_s0 .INIT=8'hE0;
  LUT3 \u_usb_device_controller/rxdat_o_d_1_s0  (
    .F(u_usb_device_controller_rxdat_o_d[1]),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_rxdat_d2[1]) 
);
defparam \u_usb_device_controller/rxdat_o_d_1_s0 .INIT=8'hE0;
  LUT3 \u_usb_device_controller/rxdat_o_d_2_s0  (
    .F(u_usb_device_controller_rxdat_o_d[2]),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_rxdat_d2[2]) 
);
defparam \u_usb_device_controller/rxdat_o_d_2_s0 .INIT=8'hE0;
  LUT3 \u_usb_device_controller/rxdat_o_d_3_s0  (
    .F(u_usb_device_controller_rxdat_o_d[3]),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_rxdat_d2[3]) 
);
defparam \u_usb_device_controller/rxdat_o_d_3_s0 .INIT=8'hE0;
  LUT3 \u_usb_device_controller/rxdat_o_d_4_s0  (
    .F(u_usb_device_controller_rxdat_o_d[4]),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_rxdat_d2[4]) 
);
defparam \u_usb_device_controller/rxdat_o_d_4_s0 .INIT=8'hE0;
  LUT3 \u_usb_device_controller/rxdat_o_d_5_s0  (
    .F(u_usb_device_controller_rxdat_o_d[5]),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_rxdat_d2[5]) 
);
defparam \u_usb_device_controller/rxdat_o_d_5_s0 .INIT=8'hE0;
  LUT3 \u_usb_device_controller/rxdat_o_d_6_s0  (
    .F(u_usb_device_controller_rxdat_o_d[6]),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_rxdat_d2[6]) 
);
defparam \u_usb_device_controller/rxdat_o_d_6_s0 .INIT=8'hE0;
  LUT3 \u_usb_device_controller/rxdat_o_d_7_s0  (
    .F(u_usb_device_controller_rxdat_o_d[7]),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_rxdat_d2[7]) 
);
defparam \u_usb_device_controller/rxdat_o_d_7_s0 .INIT=8'hE0;
  LUT3 \u_usb_device_controller/n2393_s3  (
    .F(u_usb_device_controller_n2393),
    .I0(u_usb_device_controller_rxact_o_d),
    .I1(u_usb_device_controller_setup_o_d),
    .I2(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n2393_s3 .INIT=8'hE0;
  LUT4 \u_usb_device_controller/n1595_s17  (
    .F(u_usb_device_controller_n1595),
    .I0(u_usb_device_controller_n1585),
    .I1(u_usb_device_controller_n1615_15),
    .I2(u_usb_device_controller_s_bufptr[10]),
    .I3(u_usb_device_controller_n1595_23) 
);
defparam \u_usb_device_controller/n1595_s17 .INIT=16'h0EE0;
  LUT4 \u_usb_device_controller/n1601_s17  (
    .F(u_usb_device_controller_n1601),
    .I0(u_usb_device_controller_n1585),
    .I1(u_usb_device_controller_n1615_15),
    .I2(u_usb_device_controller_s_bufptr[7]),
    .I3(u_usb_device_controller_n1601_23) 
);
defparam \u_usb_device_controller/n1601_s17 .INIT=16'h0EE0;
  LUT4 \u_usb_device_controller/n1607_s17  (
    .F(u_usb_device_controller_n1607),
    .I0(u_usb_device_controller_n1585),
    .I1(u_usb_device_controller_n1615_15),
    .I2(u_usb_device_controller_s_bufptr[4]),
    .I3(u_usb_device_controller_n1607_23) 
);
defparam \u_usb_device_controller/n1607_s17 .INIT=16'h0EE0;
  LUT4 \u_usb_device_controller/n1613_s16  (
    .F(u_usb_device_controller_n1613),
    .I0(u_usb_device_controller_n1585),
    .I1(u_usb_device_controller_n1615_15),
    .I2(u_usb_device_controller_s_bufptr[0]),
    .I3(u_usb_device_controller_s_bufptr[1]) 
);
defparam \u_usb_device_controller/n1613_s16 .INIT=16'h0EE0;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s23  (
    .F(u_usb_device_controller_u_usb_packet_n328_29),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid[0]),
    .I1(u_usb_device_controller_usb_transact_inst_n1080_53),
    .I2(u_usb_device_controller_usb_transact_inst_n1072_18),
    .I3(u_usb_device_controller_usb_transact_inst_n1157_28) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s23 .INIT=16'h1410;
  LUT4 \u_usb_device_controller/u_usb_packet/n328_s24  (
    .F(u_usb_device_controller_u_usb_packet_n328_31),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid[1]),
    .I1(u_usb_device_controller_usb_transact_inst_n1080_53),
    .I2(u_usb_device_controller_usb_transact_inst_n1072_18),
    .I3(u_usb_device_controller_usb_transact_inst_n1157_28) 
);
defparam \u_usb_device_controller/u_usb_packet/n328_s24 .INIT=16'h1410;
  LUT4 \u_usb_device_controller/usbc_dsclen_1_s18  (
    .F(u_usb_device_controller_usbc_dsclen_1_24),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscinx[3]),
    .I1(u_usb_device_controller_usb_control_inst_n1836_11),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s18 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usbc_dsclen_1_s19  (
    .F(u_usb_device_controller_usbc_dsclen_1_26),
    .I0(desc_strvendor_len_i_d[1]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscinx[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscinx[2]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscinx[0]) 
);
defparam \u_usb_device_controller/usbc_dsclen_1_s19 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/usbc_dsclen_0_s21  (
    .F(u_usb_device_controller_usbc_dsclen_0_28),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dsctyp[0]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dsctyp[1]),
    .I2(u_usb_device_controller_usb_control_inst_n1836_10),
    .I3(u_usb_device_controller_usbc_dsclen_0_17) 
);
defparam \u_usb_device_controller/usbc_dsclen_0_s21 .INIT=16'h00BF;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1068_s11  (
    .F(u_usb_device_controller_usb_transact_inst_n1068_18),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_usb_transact_inst_n1565_7),
    .I2(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I3(u_usb_device_controller_u_usb_packet_s_rxvalid) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1068_s11 .INIT=16'h7000;
  LUT4 \u_usb_device_controller/u_usb_packet/crc16_buf_15_s7  (
    .F(u_usb_device_controller_u_usb_packet_crc16_buf_15_14),
    .I0(u_usb_device_controller_u_usb_packet_s_rxerror),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I2(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I3(u_usb_device_controller_u_usb_packet_n912_14) 
);
defparam \u_usb_device_controller/u_usb_packet/crc16_buf_15_s7 .INIT=16'h4000;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1086_s45  (
    .F(u_usb_device_controller_usb_transact_inst_n1086_52),
    .I0(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I1(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I2(u_usb_device_controller_usb_transact_inst_n1064_16) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1086_s45 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1111_s16  (
    .F(u_usb_device_controller_usb_transact_inst_n1111_22),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I1(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I2(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I3(u_usb_device_controller_u_usb_packet_s_rxvalid) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1111_s16 .INIT=16'h4000;
  LUT3 \u_usb_device_controller/usb_transact_inst/s_endpt_0_s5  (
    .F(u_usb_device_controller_usb_transact_inst_s_endpt_0_9),
    .I0(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I1(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I2(u_usb_device_controller_usb_transact_inst_s_endpt_0_7) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_endpt_0_s5 .INIT=8'h80;
  LUT3 \u_usb_device_controller/n2393_s4  (
    .F(u_usb_device_controller_n2393_9),
    .I0(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I1(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I2(u_usb_device_controller_usb_transact_inst_n1095_45) 
);
defparam \u_usb_device_controller/n2393_s4 .INIT=8'h80;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_endpt_3_s3  (
    .F(u_usb_device_controller_usb_transact_inst_s_endpt_3),
    .I0(u_usb_device_controller_usb_transact_inst_s_sof),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I2(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I3(u_usb_device_controller_usb_transact_inst_n1041) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_endpt_3_s3 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/u_usb_packet/n773_s3  (
    .F(u_usb_device_controller_u_usb_packet_n773),
    .I0(u_usb_device_controller_u_usb_packet_n774_6),
    .I1(u_usb_device_controller_u_usb_packet_n912_10),
    .I2(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n773_s3 .INIT=16'hFFF6;
  LUT4 \u_usb_device_controller/u_usb_packet/n769_s3  (
    .F(u_usb_device_controller_u_usb_packet_n769),
    .I0(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I1(u_usb_device_controller_u_usb_packet_crc16_buf_15_12),
    .I2(u_usb_device_controller_u_usb_packet_n912_9),
    .I3(u_usb_device_controller_u_usb_packet_n770_6) 
);
defparam \u_usb_device_controller/u_usb_packet/n769_s3 .INIT=16'hEFFE;
  LUT4 \u_usb_device_controller/u_usb_packet/n772_s3  (
    .F(u_usb_device_controller_u_usb_packet_n772),
    .I0(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I1(u_usb_device_controller_u_usb_packet_crc16_buf_15_12),
    .I2(u_usb_device_controller_u_usb_packet_n912_10),
    .I3(u_usb_device_controller_u_usb_packet_n771_6) 
);
defparam \u_usb_device_controller/u_usb_packet/n772_s3 .INIT=16'hEFFE;
  LUT3 \u_usb_device_controller/u_usb_packet/n762_s2  (
    .F(u_usb_device_controller_u_usb_packet_n762),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[6]),
    .I1(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n762_s2 .INIT=8'hFE;
  LUT3 \u_usb_device_controller/u_usb_packet/n763_s2  (
    .F(u_usb_device_controller_u_usb_packet_n763),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[5]),
    .I1(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n763_s2 .INIT=8'hFE;
  LUT3 \u_usb_device_controller/u_usb_packet/n765_s2  (
    .F(u_usb_device_controller_u_usb_packet_n765),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[3]),
    .I1(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n765_s2 .INIT=8'hFE;
  LUT3 \u_usb_device_controller/u_usb_packet/n766_s2  (
    .F(u_usb_device_controller_u_usb_packet_n766),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[2]),
    .I1(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I2(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n766_s2 .INIT=8'hFE;
  LUT4 \u_usb_device_controller/u_usb_packet/n767_s8  (
    .F(u_usb_device_controller_u_usb_packet_n767),
    .I0(u_usb_device_controller_u_usb_packet_crc16_buf[1]),
    .I1(u_usb_device_controller_u_usb_packet_n767_6),
    .I2(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n767_s8 .INIT=16'hFFF9;
  LUT4 \u_usb_device_controller/u_usb_packet/n770_s7  (
    .F(u_usb_device_controller_u_usb_packet_n770),
    .I0(u_usb_device_controller_u_usb_packet_n770_6),
    .I1(u_usb_device_controller_u_usb_packet_n771_7),
    .I2(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n770_s7 .INIT=16'hFFF6;
  LUT4 \u_usb_device_controller/u_usb_packet/n771_s13  (
    .F(u_usb_device_controller_u_usb_packet_n771),
    .I0(u_usb_device_controller_u_usb_packet_n771_6),
    .I1(u_usb_device_controller_u_usb_packet_n771_7),
    .I2(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n771_s13 .INIT=16'hFFF6;
  LUT4 \u_usb_device_controller/u_usb_packet/n774_s8  (
    .F(u_usb_device_controller_u_usb_packet_n774),
    .I0(u_usb_device_controller_u_usb_packet_n774_6),
    .I1(u_usb_device_controller_u_usb_packet_n774_7),
    .I2(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I3(u_usb_device_controller_u_usb_packet_crc16_buf_15_12) 
);
defparam \u_usb_device_controller/u_usb_packet/n774_s8 .INIT=16'hFFF6;
  LUT4 \u_usb_device_controller/u_usb_packet/n784_s14  (
    .F(u_usb_device_controller_u_usb_packet_n784_20),
    .I0(u_usb_device_controller_u_usb_packet_n626_42),
    .I1(u_usb_device_controller_usb_transact_inst_n1072_18),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[5]),
    .I3(u_usb_device_controller_usb_transact_inst_n1091_50) 
);
defparam \u_usb_device_controller/u_usb_packet/n784_s14 .INIT=16'h0015;
  LUT4 \u_usb_device_controller/u_usb_init/s_state_2_s14  (
    .F(u_usb_device_controller_u_usb_init_s_state_2),
    .I0(u_usb_device_controller_u_usb_init_n212_29),
    .I1(u_usb_device_controller_u_usb_init_s_state[3]),
    .I2(u_usb_device_controller_u_usb_init_s_state[2]),
    .I3(u_usb_device_controller_u_usb_init_s_state_2_14) 
);
defparam \u_usb_device_controller/u_usb_init/s_state_2_s14 .INIT=16'hEF00;
  LUT4 \u_usb_device_controller/usb_control_inst/n1652_s18  (
    .F(u_usb_device_controller_usb_control_inst_n1652_24),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscoff[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_dscoff[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_dscoff[0]),
    .I3(u_usb_device_controller_usb_control_inst_usbc_dscoff[1]) 
);
defparam \u_usb_device_controller/usb_control_inst/n1652_s18 .INIT=16'h8000;
  LUT4 \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s15  (
    .F(u_usb_device_controller_usb_control_inst_s_sendbyte_7),
    .I0(u_usb_device_controller_usb_control_inst_s_sendbyte_7_15),
    .I1(u_usb_device_controller_usb_control_inst_s_state[6]),
    .I2(u_usb_device_controller_usb_control_inst_s_answerptr_5_14),
    .I3(u_usb_device_controller_usb_control_inst_s_sendbyte_7_13) 
);
defparam \u_usb_device_controller/usb_control_inst/s_sendbyte_7_s15 .INIT=16'hBF00;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1091_s49  (
    .F(u_usb_device_controller_usb_transact_inst_n1091_56),
    .I0(u_usb_device_controller_usb_transact_inst_n1091_54),
    .I1(u_usb_device_controller_u_usb_packet_n800_6),
    .I2(u_usb_device_controller_usb_transact_inst_n1091_50),
    .I3(u_usb_device_controller_u_usb_packet_n626_42) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1091_s49 .INIT=16'hFFE0;
  LUT3 \u_usb_device_controller/usb_transact_inst/n1140_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1140),
    .I0(u_usb_device_controller_u_usb_init_highspeed_o_d),
    .I1(u_usb_device_controller_usb_transact_inst_n1142_25),
    .I2(u_usb_device_controller_usb_transact_inst_n1140_22) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1140_s19 .INIT=8'hF1;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s15  (
    .F(u_usb_device_controller_usb_transact_inst_s_sendpid_3_23),
    .I0(u_usb_device_controller_usb_transact_inst_n1099_49),
    .I1(u_usb_device_controller_usb_transact_inst_s_ping),
    .I2(u_usb_device_controller_usb_transact_inst_s_in),
    .I3(u_usb_device_controller_usb_transact_inst_n1163_24) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_sendpid_3_s15 .INIT=16'h0155;
  LUT4 \u_usb_device_controller/u_usb_packet/n622_s41  (
    .F(u_usb_device_controller_u_usb_packet_n622),
    .I0(u_usb_device_controller_u_usb_packet_n784_20),
    .I1(u_usb_device_controller_u_usb_packet_s_txfirst),
    .I2(u_usb_device_controller_u_usb_packet_s_txready),
    .I3(u_usb_device_controller_u_usb_packet_n615_49) 
);
defparam \u_usb_device_controller/u_usb_packet/n622_s41 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1107_s43  (
    .F(u_usb_device_controller_usb_transact_inst_n1107_48),
    .I0(u_usb_device_controller_usb_transact_inst_n1068_18),
    .I1(u_usb_device_controller_usb_transact_inst_n1088_48),
    .I2(u_usb_device_controller_usb_transact_inst_n1111),
    .I3(u_usb_device_controller_usb_transact_inst_n1064_23) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1107_s43 .INIT=16'hF800;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1064_s18  (
    .F(u_usb_device_controller_usb_transact_inst_n1064_25),
    .I0(u_usb_device_controller_usb_transact_inst_n1068_16),
    .I1(u_usb_device_controller_usb_transact_inst_n1068_18),
    .I2(u_usb_device_controller_usb_transact_inst_n1088_48),
    .I3(u_usb_device_controller_usb_transact_inst_s_in) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1064_s18 .INIT=16'h1500;
  LUT4 \u_usb_device_controller/usb_transact_inst/s_endpt_0_s6  (
    .F(u_usb_device_controller_usb_transact_inst_s_endpt_0),
    .I0(u_usb_device_controller_usb_transact_inst_s_sof),
    .I1(u_usb_device_controller_u_usb_packet_usbp_rxact),
    .I2(u_usb_device_controller_u_usb_packet_s_rxvalid),
    .I3(u_usb_device_controller_usb_transact_inst_s_endpt_0_7) 
);
defparam \u_usb_device_controller/usb_transact_inst/s_endpt_0_s6 .INIT=16'h4000;
  LUT4 \u_usb_device_controller/usb_control_inst/n1674_s38  (
    .F(u_usb_device_controller_usb_control_inst_n1674_44),
    .I0(u_usb_device_controller_usb_control_inst_n1680_50),
    .I1(u_usb_device_controller_usb_control_inst_n1474_3),
    .I2(u_usb_device_controller_usb_control_inst_n1483_3),
    .I3(u_usb_device_controller_usb_transact_inst_txpop_o_d_5) 
);
defparam \u_usb_device_controller/usb_control_inst/n1674_s38 .INIT=16'hBF00;
  LUT3 \u_usb_device_controller/usb_control_inst/s_ctlparam_7_s6  (
    .F(u_usb_device_controller_usb_control_inst_s_ctlparam_7),
    .I0(u_usb_device_controller_u_usb_init_utmi_reset_o_d),
    .I1(u_usb_device_controller_usb_control_inst_n1836_15),
    .I2(u_usb_device_controller_usb_control_inst_s_ctlparam_7_7) 
);
defparam \u_usb_device_controller/usb_control_inst/s_ctlparam_7_s6 .INIT=8'h40;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1099_s45  (
    .F(u_usb_device_controller_usb_transact_inst_n1099),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I3(u_usb_device_controller_usb_transact_inst_n1099_47) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1099_s45 .INIT=16'h20FF;
  LUT4 \u_usb_device_controller/usb_transact_inst/wait_count_9_s4  (
    .F(u_usb_device_controller_usb_transact_inst_wait_count_9),
    .I0(u_usb_device_controller_usb_transact_inst_s_sendpid_3),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[4]),
    .I2(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_41) 
);
defparam \u_usb_device_controller/usb_transact_inst/wait_count_9_s4 .INIT=16'hDF00;
  LUT4 \u_usb_device_controller/s_bufptr_1_s4  (
    .F(u_usb_device_controller_s_bufptr_1),
    .I0(u_usb_device_controller_usb_transact_inst_txpop_o_d_9),
    .I1(u_usb_device_controller_usb_transact_inst_txpop_o_d_5),
    .I2(u_usb_device_controller_n1615_15),
    .I3(u_usb_device_controller_n1593_24) 
);
defparam \u_usb_device_controller/s_bufptr_1_s4 .INIT=16'h4F00;
  LUT3 \u_usb_device_controller/usb_control_inst/usbc_dscrd_s1  (
    .F(u_usb_device_controller_usb_control_inst_usbc_dscrd),
    .I0(u_usb_device_controller_usb_control_inst_usbc_dscrd_4),
    .I1(u_usb_device_controller_usb_transact_inst_txpop_o_d_9),
    .I2(u_usb_device_controller_usb_transact_inst_txpop_o_d_5) 
);
defparam \u_usb_device_controller/usb_control_inst/usbc_dscrd_s1 .INIT=8'hBA;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1064_s19  (
    .F(u_usb_device_controller_usb_transact_inst_n1064_27),
    .I0(u_usb_device_controller_usb_transact_inst_n1080_53),
    .I1(u_usb_device_controller_usb_transact_inst_s_state[8]),
    .I2(u_usb_device_controller_usb_transact_inst_s_state[9]),
    .I3(u_usb_device_controller_usb_transact_inst_n1157_28) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1064_s19 .INIT=16'h0200;
  LUT4 \u_usb_device_controller/usb_transact_inst/n1138_s33  (
    .F(u_usb_device_controller_usb_transact_inst_n1138_43),
    .I0(u_usb_device_controller_usb_transact_inst_n1157_23),
    .I1(u_usb_device_controller_usb_transact_inst_n1064_16),
    .I2(u_usb_device_controller_usb_transact_inst_n1138_24),
    .I3(u_usb_device_controller_usb_transact_inst_n1138_37) 
);
defparam \u_usb_device_controller/usb_transact_inst/n1138_s33 .INIT=16'h00FE;
  LUT4 \u_usb_device_controller/n1716_s2  (
    .F(u_usb_device_controller_n1716),
    .I0(u_usb_device_controller_rxval_d0),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1716_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1714_s2  (
    .F(u_usb_device_controller_n1714),
    .I0(u_usb_device_controller_rxdat_d0[0]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1714_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1713_s2  (
    .F(u_usb_device_controller_n1713),
    .I0(u_usb_device_controller_rxdat_d0[1]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1713_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1712_s2  (
    .F(u_usb_device_controller_n1712),
    .I0(u_usb_device_controller_rxdat_d0[2]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1712_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1711_s2  (
    .F(u_usb_device_controller_n1711),
    .I0(u_usb_device_controller_rxdat_d0[3]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1711_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1710_s2  (
    .F(u_usb_device_controller_n1710),
    .I0(u_usb_device_controller_rxdat_d0[4]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1710_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1709_s2  (
    .F(u_usb_device_controller_n1709),
    .I0(u_usb_device_controller_rxdat_d0[5]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1709_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1708_s2  (
    .F(u_usb_device_controller_n1708),
    .I0(u_usb_device_controller_rxdat_d0[6]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1708_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1707_s2  (
    .F(u_usb_device_controller_n1707),
    .I0(u_usb_device_controller_rxdat_d0[7]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1707_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1706_s2  (
    .F(u_usb_device_controller_n1706),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[0]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1706_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1705_s2  (
    .F(u_usb_device_controller_n1705),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[1]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1705_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1704_s2  (
    .F(u_usb_device_controller_n1704),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[2]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1704_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1703_s2  (
    .F(u_usb_device_controller_n1703),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[3]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1703_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1702_s2  (
    .F(u_usb_device_controller_n1702),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[4]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1702_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1701_s2  (
    .F(u_usb_device_controller_n1701),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[5]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1701_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1700_s2  (
    .F(u_usb_device_controller_n1700),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[6]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1700_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1699_s2  (
    .F(u_usb_device_controller_n1699),
    .I0(u_usb_device_controller_u_usb_packet_usbt_rxdat[7]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1699_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1760_s2  (
    .F(u_usb_device_controller_n1760),
    .I0(u_usb_device_controller_rxdat_d1[7]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1760_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1761_s2  (
    .F(u_usb_device_controller_n1761),
    .I0(u_usb_device_controller_rxdat_d1[6]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1761_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1762_s2  (
    .F(u_usb_device_controller_n1762),
    .I0(u_usb_device_controller_rxdat_d1[5]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1762_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1763_s2  (
    .F(u_usb_device_controller_n1763),
    .I0(u_usb_device_controller_rxdat_d1[4]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1763_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1764_s2  (
    .F(u_usb_device_controller_n1764),
    .I0(u_usb_device_controller_rxdat_d1[3]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1764_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1765_s2  (
    .F(u_usb_device_controller_n1765),
    .I0(u_usb_device_controller_rxdat_d1[2]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1765_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1766_s2  (
    .F(u_usb_device_controller_n1766),
    .I0(u_usb_device_controller_rxdat_d1[1]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1766_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1767_s2  (
    .F(u_usb_device_controller_n1767),
    .I0(u_usb_device_controller_rxdat_d1[0]),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1767_s2 .INIT=16'hA800;
  LUT4 \u_usb_device_controller/n1770_s2  (
    .F(u_usb_device_controller_n1770),
    .I0(u_usb_device_controller_rxval_d1),
    .I1(u_usb_device_controller_rxact_o_d),
    .I2(u_usb_device_controller_setup_o_d),
    .I3(u_usb_device_controller_n2393_9) 
);
defparam \u_usb_device_controller/n1770_s2 .INIT=16'hA800;
  DFFR \u_usb_device_controller/u_usb_init/s_timer1_0_s1  (
    .Q(u_usb_device_controller_u_usb_init_s_timer1[0]),
    .D(u_usb_device_controller_u_usb_init_n241),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_u_usb_init_n242) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer1_0_s1 .INIT=1'b0;
  DFFR \u_usb_device_controller/u_usb_init/s_timer2_0_s1  (
    .Q(u_usb_device_controller_u_usb_init_s_timer2[0]),
    .D(u_usb_device_controller_u_usb_init_n279),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_u_usb_init_n280) 
);
defparam \u_usb_device_controller/u_usb_init/s_timer2_0_s1 .INIT=1'b0;
  DFF \u_usb_device_controller/usb_control_inst/s_setupptr_0_s5  (
    .Q(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .D(u_usb_device_controller_usb_control_inst_n1699_15),
    .CLK(clk_i_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_setupptr_0_s5 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_1_s4  (
    .Q(u_usb_device_controller_halt_out[1]),
    .D(u_usb_device_controller_n340),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_1_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_2_s4  (
    .Q(u_usb_device_controller_halt_in[2]),
    .D(u_usb_device_controller_n395),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_2_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_2_s4  (
    .Q(u_usb_device_controller_halt_out[2]),
    .D(u_usb_device_controller_n398),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_2_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_3_s4  (
    .Q(u_usb_device_controller_halt_in[3]),
    .D(u_usb_device_controller_n453),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_3_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_3_s4  (
    .Q(u_usb_device_controller_halt_out[3]),
    .D(u_usb_device_controller_n456),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_3_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_4_s4  (
    .Q(u_usb_device_controller_halt_in[4]),
    .D(u_usb_device_controller_n513),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_4_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_4_s4  (
    .Q(u_usb_device_controller_halt_out[4]),
    .D(u_usb_device_controller_n516),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_4_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_5_s4  (
    .Q(u_usb_device_controller_halt_in[5]),
    .D(u_usb_device_controller_n571),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_5_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_5_s4  (
    .Q(u_usb_device_controller_halt_out[5]),
    .D(u_usb_device_controller_n574),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_5_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_6_s4  (
    .Q(u_usb_device_controller_halt_in[6]),
    .D(u_usb_device_controller_n631),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_6_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_6_s4  (
    .Q(u_usb_device_controller_halt_out[6]),
    .D(u_usb_device_controller_n634),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_6_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_7_s4  (
    .Q(u_usb_device_controller_halt_in[7]),
    .D(u_usb_device_controller_n691),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_7_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_7_s4  (
    .Q(u_usb_device_controller_halt_out[7]),
    .D(u_usb_device_controller_n694),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_7_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_8_s4  (
    .Q(u_usb_device_controller_halt_in[8]),
    .D(u_usb_device_controller_n753),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_8_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_8_s4  (
    .Q(u_usb_device_controller_halt_out[8]),
    .D(u_usb_device_controller_n756),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_8_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_9_s4  (
    .Q(u_usb_device_controller_halt_in[9]),
    .D(u_usb_device_controller_n811),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_9_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_9_s4  (
    .Q(u_usb_device_controller_halt_out[9]),
    .D(u_usb_device_controller_n814),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_9_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_10_s4  (
    .Q(u_usb_device_controller_halt_in[10]),
    .D(u_usb_device_controller_n871),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_10_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_10_s4  (
    .Q(u_usb_device_controller_halt_out[10]),
    .D(u_usb_device_controller_n874),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_10_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_11_s4  (
    .Q(u_usb_device_controller_halt_in[11]),
    .D(u_usb_device_controller_n931),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_11_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_11_s4  (
    .Q(u_usb_device_controller_halt_out[11]),
    .D(u_usb_device_controller_n934),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_11_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_12_s4  (
    .Q(u_usb_device_controller_halt_in[12]),
    .D(u_usb_device_controller_n993),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_12_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_12_s4  (
    .Q(u_usb_device_controller_halt_out[12]),
    .D(u_usb_device_controller_n996),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_12_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_13_s4  (
    .Q(u_usb_device_controller_halt_in[13]),
    .D(u_usb_device_controller_n1053),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_13_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_13_s4  (
    .Q(u_usb_device_controller_halt_out[13]),
    .D(u_usb_device_controller_n1056),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_13_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_14_s4  (
    .Q(u_usb_device_controller_halt_in[14]),
    .D(u_usb_device_controller_n1115),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_14_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_14_s4  (
    .Q(u_usb_device_controller_halt_out[14]),
    .D(u_usb_device_controller_n1118),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_14_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_15_s4  (
    .Q(u_usb_device_controller_halt_in[15]),
    .D(u_usb_device_controller_n1177),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_15_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_out_15_s4  (
    .Q(u_usb_device_controller_halt_out[15]),
    .D(u_usb_device_controller_n1180),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_out_15_s4 .INIT=1'b0;
  DFFR \u_usb_device_controller/halt_in_1_s4  (
    .Q(u_usb_device_controller_halt_in[1]),
    .D(u_usb_device_controller_n337),
    .CLK(clk_i_d),
    .RESET(u_usb_device_controller_n2219) 
);
defparam \u_usb_device_controller/halt_in_1_s4 .INIT=1'b0;
  LUT2 \u_usb_device_controller/u_usb_init/n241_s3  (
    .F(u_usb_device_controller_u_usb_init_n241),
    .I0(u_usb_device_controller_u_usb_init_s_timer1[0]),
    .I1(reset_i_d) 
);
defparam \u_usb_device_controller/u_usb_init/n241_s3 .INIT=4'h9;
  LUT2 \u_usb_device_controller/u_usb_init/n279_s3  (
    .F(u_usb_device_controller_u_usb_init_n279),
    .I0(reset_i_d),
    .I1(u_usb_device_controller_u_usb_init_s_timer2[0]) 
);
defparam \u_usb_device_controller/u_usb_init/n279_s3 .INIT=4'h9;
  LUT4 \u_usb_device_controller/usb_control_inst/n1699_s10  (
    .F(u_usb_device_controller_usb_control_inst_n1699_15),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I1(u_usb_device_controller_usb_control_inst_n1836_15),
    .I2(u_usb_device_controller_usb_control_inst_s_setupptr_2_12),
    .I3(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/n1699_s10 .INIT=16'hAA46;
  LUT2 \u_usb_device_controller/usb_control_inst/n1699_s11  (
    .F(u_usb_device_controller_usb_control_inst_n1699),
    .I0(u_usb_device_controller_usb_control_inst_s_setupptr[0]),
    .I1(u_usb_device_controller_usb_control_inst_n1836_15) 
);
defparam \u_usb_device_controller/usb_control_inst/n1699_s11 .INIT=4'h4;
  LUT3 \u_usb_device_controller/usb_control_inst/s_setupptr_2_s8  (
    .F(u_usb_device_controller_usb_control_inst_s_setupptr_2),
    .I0(u_usb_device_controller_usb_control_inst_n1836_15),
    .I1(u_usb_device_controller_usb_control_inst_s_setupptr_2_12),
    .I2(u_usb_device_controller_u_usb_init_utmi_reset_o_d) 
);
defparam \u_usb_device_controller/usb_control_inst/s_setupptr_2_s8 .INIT=8'h0E;
  LUT3 \u_usb_device_controller/n340_s5  (
    .F(u_usb_device_controller_n340),
    .I0(u_usb_device_controller_halt_out[1]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[1]) 
);
defparam \u_usb_device_controller/n340_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n395_s5  (
    .F(u_usb_device_controller_n395),
    .I0(u_usb_device_controller_halt_in[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[2]) 
);
defparam \u_usb_device_controller/n395_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n398_s5  (
    .F(u_usb_device_controller_n398),
    .I0(u_usb_device_controller_halt_out[2]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[2]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[2]) 
);
defparam \u_usb_device_controller/n398_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n453_s5  (
    .F(u_usb_device_controller_n453),
    .I0(u_usb_device_controller_halt_in[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[3]) 
);
defparam \u_usb_device_controller/n453_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n456_s5  (
    .F(u_usb_device_controller_n456),
    .I0(u_usb_device_controller_halt_out[3]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[3]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[3]) 
);
defparam \u_usb_device_controller/n456_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n513_s5  (
    .F(u_usb_device_controller_n513),
    .I0(u_usb_device_controller_halt_in[4]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[4]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[4]) 
);
defparam \u_usb_device_controller/n513_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n516_s5  (
    .F(u_usb_device_controller_n516),
    .I0(u_usb_device_controller_halt_out[4]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[4]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[4]) 
);
defparam \u_usb_device_controller/n516_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n571_s5  (
    .F(u_usb_device_controller_n571),
    .I0(u_usb_device_controller_halt_in[5]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[5]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[5]) 
);
defparam \u_usb_device_controller/n571_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n574_s5  (
    .F(u_usb_device_controller_n574),
    .I0(u_usb_device_controller_halt_out[5]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[5]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[5]) 
);
defparam \u_usb_device_controller/n574_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n631_s5  (
    .F(u_usb_device_controller_n631),
    .I0(u_usb_device_controller_halt_in[6]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[6]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[6]) 
);
defparam \u_usb_device_controller/n631_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n634_s5  (
    .F(u_usb_device_controller_n634),
    .I0(u_usb_device_controller_halt_out[6]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[6]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[6]) 
);
defparam \u_usb_device_controller/n634_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n691_s5  (
    .F(u_usb_device_controller_n691),
    .I0(u_usb_device_controller_halt_in[7]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[7]) 
);
defparam \u_usb_device_controller/n691_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n694_s5  (
    .F(u_usb_device_controller_n694),
    .I0(u_usb_device_controller_halt_out[7]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[7]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[7]) 
);
defparam \u_usb_device_controller/n694_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n753_s5  (
    .F(u_usb_device_controller_n753),
    .I0(u_usb_device_controller_halt_in[8]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[8]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[8]) 
);
defparam \u_usb_device_controller/n753_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n756_s5  (
    .F(u_usb_device_controller_n756),
    .I0(u_usb_device_controller_halt_out[8]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[8]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[8]) 
);
defparam \u_usb_device_controller/n756_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n811_s5  (
    .F(u_usb_device_controller_n811),
    .I0(u_usb_device_controller_halt_in[9]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[9]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[9]) 
);
defparam \u_usb_device_controller/n811_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n814_s5  (
    .F(u_usb_device_controller_n814),
    .I0(u_usb_device_controller_halt_out[9]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[9]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[9]) 
);
defparam \u_usb_device_controller/n814_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n871_s5  (
    .F(u_usb_device_controller_n871),
    .I0(u_usb_device_controller_halt_in[10]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[10]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[10]) 
);
defparam \u_usb_device_controller/n871_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n874_s5  (
    .F(u_usb_device_controller_n874),
    .I0(u_usb_device_controller_halt_out[10]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[10]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[10]) 
);
defparam \u_usb_device_controller/n874_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n931_s5  (
    .F(u_usb_device_controller_n931),
    .I0(u_usb_device_controller_halt_in[11]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[11]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[11]) 
);
defparam \u_usb_device_controller/n931_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n934_s5  (
    .F(u_usb_device_controller_n934),
    .I0(u_usb_device_controller_halt_out[11]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[11]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[11]) 
);
defparam \u_usb_device_controller/n934_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n993_s5  (
    .F(u_usb_device_controller_n993),
    .I0(u_usb_device_controller_halt_in[12]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[12]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[12]) 
);
defparam \u_usb_device_controller/n993_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n996_s5  (
    .F(u_usb_device_controller_n996),
    .I0(u_usb_device_controller_halt_out[12]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[12]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[12]) 
);
defparam \u_usb_device_controller/n996_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n1053_s5  (
    .F(u_usb_device_controller_n1053),
    .I0(u_usb_device_controller_halt_in[13]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[13]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[13]) 
);
defparam \u_usb_device_controller/n1053_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n1056_s5  (
    .F(u_usb_device_controller_n1056),
    .I0(u_usb_device_controller_halt_out[13]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[13]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[13]) 
);
defparam \u_usb_device_controller/n1056_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n1115_s5  (
    .F(u_usb_device_controller_n1115),
    .I0(u_usb_device_controller_halt_in[14]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[14]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[14]) 
);
defparam \u_usb_device_controller/n1115_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n1118_s5  (
    .F(u_usb_device_controller_n1118),
    .I0(u_usb_device_controller_halt_out[14]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[14]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[14]) 
);
defparam \u_usb_device_controller/n1118_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n1177_s5  (
    .F(u_usb_device_controller_n1177),
    .I0(u_usb_device_controller_halt_in[15]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[15]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[15]) 
);
defparam \u_usb_device_controller/n1177_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n1180_s5  (
    .F(u_usb_device_controller_n1180),
    .I0(u_usb_device_controller_halt_out[15]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_out[15]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_out[15]) 
);
defparam \u_usb_device_controller/n1180_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n337_s5  (
    .F(u_usb_device_controller_n337),
    .I0(u_usb_device_controller_halt_in[1]),
    .I1(u_usb_device_controller_usb_control_inst_usbc_clr_in[1]),
    .I2(u_usb_device_controller_usb_control_inst_usbc_sethlt_in[1]) 
);
defparam \u_usb_device_controller/n337_s5 .INIT=8'h32;
  LUT3 \u_usb_device_controller/n2024_s5  (
    .F(u_usb_device_controller_n2024),
    .I0(u_usb_device_controller_n2024_11),
    .I1(desc_oscfg_addr_i_d[9]),
    .I2(u_usb_device_controller_n2024_4) 
);
defparam \u_usb_device_controller/n2024_s5 .INIT=8'hCA;
  LUT3 \u_usb_device_controller/n2024_s6  (
    .F(u_usb_device_controller_n2024_11),
    .I0(u_usb_device_controller_descrom_start_9),
    .I1(GND),
    .I2(u_usb_device_controller_n2015_2) 
);
defparam \u_usb_device_controller/n2024_s6 .INIT=8'h96;
  INV \u_usb_device_controller/u_usb_init/n316_s3  (
    .O(u_usb_device_controller_u_usb_init_n316),
    .I(reset_i_d) 
);
assign u_usb_device_controller_usb_transact_inst_T_PING_2 = u_usb_device_controller_usb_transact_inst_T_PING;
assign u_usb_device_controller_usb_transact_inst_s_setup_2 = u_usb_device_controller_usb_transact_inst_s_setup;
  GND GND_s (
    .G(GND) 
);
  VCC VCC_s (
    .V(VCC) 
);
  GSR GSR (
    .GSRI(VCC) 
);
endmodule /* USB_Device_Controller_Top */
